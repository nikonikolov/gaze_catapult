
//------> ./rtl_mgc_ioport.v 
//------------------------------------------------------------------
//                M G C _ I O P O R T _ C O M P S
//------------------------------------------------------------------

//------------------------------------------------------------------
//                       M O D U L E S
//------------------------------------------------------------------

//------------------------------------------------------------------
//-- INPUT ENTITIES
//------------------------------------------------------------------

module mgc_in_wire (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output [width-1:0] d;
  input  [width-1:0] z;

  wire   [width-1:0] d;

  assign d = z;

endmodule

//------------------------------------------------------------------

module mgc_in_wire_en (ld, d, lz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output [width-1:0] d;
  output             lz;
  input  [width-1:0] z;

  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;

endmodule

//------------------------------------------------------------------

module mgc_in_wire_wait (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;

  wire               vd;
  wire   [width-1:0] d;
  wire               lz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;

endmodule
//------------------------------------------------------------------

module mgc_chan_in (ld, vd, d, lz, vz, z, size, req_size, sizez, sizelz);

  parameter integer rscid = 1;
  parameter integer width = 8;
  parameter integer sz_width = 8;

  input              ld;
  output             vd;
  output [width-1:0] d;
  output             lz;
  input              vz;
  input  [width-1:0] z;
  output [sz_width-1:0] size;
  input              req_size;
  input  [sz_width-1:0] sizez;
  output             sizelz;


  wire               vd;
  wire   [width-1:0] d;
  wire               lz;
  wire   [sz_width-1:0] size;
  wire               sizelz;

  assign d = z;
  assign lz = ld;
  assign vd = vz;
  assign size = sizez;
  assign sizelz = req_size;

endmodule


//------------------------------------------------------------------
//-- OUTPUT ENTITIES
//------------------------------------------------------------------

module mgc_out_stdreg (d, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input    [width-1:0] d;
  output   [width-1:0] z;

  wire     [width-1:0] z;

  assign z = d;

endmodule

//------------------------------------------------------------------

module mgc_out_stdreg_en (ld, d, lz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  input  [width-1:0] d;
  output             lz;
  output [width-1:0] z;

  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;

endmodule

//------------------------------------------------------------------

module mgc_out_stdreg_wait (ld, vd, d, lz, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  input              ld;
  output             vd;
  input  [width-1:0] d;
  output             lz;
  input              vz;
  output [width-1:0] z;

  wire               vd;
  wire               lz;
  wire   [width-1:0] z;

  assign z = d;
  assign lz = ld;
  assign vd = vz;

endmodule

//------------------------------------------------------------------

module mgc_out_prereg_en (ld, d, lz, z);

    parameter integer rscid = 1;
    parameter integer width = 8;

    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;

    wire               lz;
    wire   [width-1:0] z;

    assign z = d;
    assign lz = ld;

endmodule

//------------------------------------------------------------------
//-- INOUT ENTITIES
//------------------------------------------------------------------

module mgc_inout_stdreg_en (ldin, din, ldout, dout, lzin, lzout, z);

    parameter integer rscid = 1;
    parameter integer width = 8;

    input              ldin;
    output [width-1:0] din;
    input              ldout;
    input  [width-1:0] dout;
    output             lzin;
    output             lzout;
    inout  [width-1:0] z;

    wire   [width-1:0] din;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzin = ldin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = ldout;
    assign z = ldout ? dout : {width{1'bz}};

endmodule

//------------------------------------------------------------------
module hid_tribuf( I_SIG, ENABLE, O_SIG);
  parameter integer width = 8;

  input [width-1:0] I_SIG;
  input ENABLE;
  inout [width-1:0] O_SIG;

  assign O_SIG = (ENABLE) ? I_SIG : { width{1'bz}};

endmodule
//------------------------------------------------------------------

module mgc_inout_stdreg_wait (ldin, vdin, din, ldout, vdout, dout, lzin, vzin, lzout, vzout, z);

    parameter integer rscid = 1;
    parameter integer width = 8;

    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output             lzin;
    input              vzin;
    output             lzout;
    input              vzout;
    inout  [width-1:0] z;

    wire               vdin;
    wire   [width-1:0] din;
    wire               vdout;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;
    wire   ldout_and_vzout;

    assign lzin = ldin;
    assign vdin = vzin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = ldout;
    assign vdout = vzout ;
    assign ldout_and_vzout = ldout && vzout ;

    hid_tribuf #(width) tb( .I_SIG(dout),
                            .ENABLE(ldout_and_vzout),
                            .O_SIG(z) );

endmodule

//------------------------------------------------------------------

module mgc_inout_buf_wait (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, lzin, vzin, lzout, vzout, z);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter         ph_clk  =  1'b1; // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   =  1'b1; // clock enable polarity
    parameter         ph_arst =  1'b1; // async reset polarity
    parameter         ph_srst =  1'b1; // sync reset polarity

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output             lzin;
    input              vzin;
    output             lzout;
    input              vzout;
    inout  [width-1:0] z;

    wire               lzout_buf;
    wire               vzout_buf;
    wire   [width-1:0] z_buf;
    wire               vdin;
    wire   [width-1:0] din;
    wire               vdout;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzin = ldin;
    assign vdin = vzin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = lzout_buf & ~ldin;
    assign vzout_buf = vzout & ~ldin;
    hid_tribuf #(width) tb( .I_SIG(z_buf),
                            .ENABLE((lzout_buf && (!ldin) && vzout) ),
                            .O_SIG(z)  );

    mgc_out_buf_wait
    #(
        .rscid   (rscid),
        .width   (width),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst)
    )
    BUFF
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (lzout_buf),
        .vz      (vzout_buf),
        .z       (z_buf)
    );


endmodule

module mgc_inout_fifo_wait (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, lzin, vzin, lzout, vzout, z);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer fifo_sz = 8; // fifo depth
    parameter         ph_clk  = 1'b1;  // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   = 1'b1;  // clock enable polarity
    parameter         ph_arst = 1'b1;  // async reset polarity
    parameter         ph_srst = 1'b1;  // sync reset polarity
    parameter integer ph_log2 = 3;     // log2(fifo_sz)
    parameter integer pwropt  = 0;     // pwropt

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output             lzin;
    input              vzin;
    output             lzout;
    input              vzout;
    inout  [width-1:0] z;

    wire               lzout_buf;
    wire               vzout_buf;
    wire   [width-1:0] z_buf;
    wire               comb;
    wire               vdin;
    wire   [width-1:0] din;
    wire               vdout;
    wire               lzin;
    wire               lzout;
    wire   [width-1:0] z;

    assign lzin = ldin;
    assign vdin = vzin;
    assign din = ldin ? z : {width{1'bz}};
    assign lzout = lzout_buf & ~ldin;
    assign vzout_buf = vzout & ~ldin;
    assign comb = (lzout_buf && (!ldin) && vzout);

    hid_tribuf #(width) tb2( .I_SIG(z_buf), .ENABLE(comb), .O_SIG(z)  );

    mgc_out_fifo_wait
    #(
        .rscid   (rscid),
        .width   (width),
        .fifo_sz (fifo_sz),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .ph_log2 (ph_log2),
        .pwropt  (pwropt)
    )
    FIFO
    (
        .clk   (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (lzout_buf),
        .vz      (vzout_buf),
        .z       (z_buf)
    );

endmodule

//------------------------------------------------------------------
//-- I/O SYNCHRONIZATION ENTITIES
//------------------------------------------------------------------

module mgc_io_sync (ld, lz);

    input  ld;
    output lz;

    assign lz = ld;

endmodule

module mgc_bsync_rdy (rd, rz);

    parameter integer rscid   = 0; // resource ID
    parameter ready = 1;
    parameter valid = 0;

    input  rd;
    output rz;

    wire   rz;

    assign rz = rd;

endmodule

module mgc_bsync_vld (vd, vz);

    parameter integer rscid   = 0; // resource ID
    parameter ready = 0;
    parameter valid = 1;

    output vd;
    input  vz;

    wire   vd;

    assign vd = vz;

endmodule

module mgc_bsync_rv (rd, vd, rz, vz);

    parameter integer rscid   = 0; // resource ID
    parameter ready = 1;
    parameter valid = 1;

    input  rd;
    output vd;
    output rz;
    input  vz;

    wire   vd;
    wire   rz;

    assign rz = rd;
    assign vd = vz;

endmodule

//------------------------------------------------------------------

module mgc_sync (ldin, vdin, ldout, vdout);

  input  ldin;
  output vdin;
  input  ldout;
  output vdout;

  wire   vdin;
  wire   vdout;

  assign vdin = ldout;
  assign vdout = ldin;

endmodule

///////////////////////////////////////////////////////////////////////////////
// dummy function used to preserve funccalls for modulario
// it looks like a memory read to the caller
///////////////////////////////////////////////////////////////////////////////
module funccall_inout (d, ad, bd, z, az, bz);

  parameter integer ram_id = 1;
  parameter integer width = 8;
  parameter integer addr_width = 8;

  output [width-1:0]       d;
  input  [addr_width-1:0]  ad;
  input                    bd;
  input  [width-1:0]       z;
  output [addr_width-1:0]  az;
  output                   bz;

  wire   [width-1:0]       d;
  wire   [addr_width-1:0]  az;
  wire                     bz;

  assign d  = z;
  assign az = ad;
  assign bz = bd;

endmodule


///////////////////////////////////////////////////////////////////////////////
// inlinable modular io not otherwise found in mgc_ioport
///////////////////////////////////////////////////////////////////////////////

module modulario_en_in (vd, d, vz, z);

  parameter integer rscid = 1;
  parameter integer width = 8;

  output             vd;
  output [width-1:0] d;
  input              vz;
  input  [width-1:0] z;

  wire   [width-1:0] d;
  wire               vd;

  assign d = z;
  assign vd = vz;

endmodule

//------> ./rtl_mgc_ioport_v2001.v 
//------------------------------------------------------------------

module mgc_out_reg_pos (clk, en, arst, srst, ld, d, lz, z);

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;

    reg                lz;
    reg    [width-1:0] z;

    generate
    if (ph_arst == 1'b0)
    begin: NEG_ARST
        always @(posedge clk or negedge arst)
        if (arst == 1'b0)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    else
    begin: POS_ARST
        always @(posedge clk or posedge arst)
        if (arst == 1'b1)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    endgenerate

endmodule

//------------------------------------------------------------------

module mgc_out_reg_neg (clk, en, arst, srst, ld, d, lz, z);

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;

    reg                lz;
    reg    [width-1:0] z;

    generate
    if (ph_arst == 1'b0)
    begin: NEG_ARST
        always @(negedge clk or negedge arst)
        if (arst == 1'b0)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    else
    begin: POS_ARST
        always @(negedge clk or posedge arst)
        if (arst == 1'b1)
        begin: B1
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (srst == ph_srst)
        begin: B2
            lz <= 1'b0;
            z  <= {width{1'b0}};
        end
        else if (en == ph_en)
        begin: B3
            lz <= ld;
            z  <= (ld) ? d : z;
        end
    end
    endgenerate

endmodule

//------------------------------------------------------------------

module mgc_out_reg (clk, en, arst, srst, ld, d, lz, z); // Not Supported

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_clk  =  1'b1;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    input  [width-1:0] d;
    output             lz;
    output [width-1:0] z;


    generate
    if (ph_clk == 1'b0)
    begin: NEG_EDGE

        mgc_out_reg_neg
        #(
            .rscid   (rscid),
            .width   (width),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        mgc_out_reg_neg_inst
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (ld),
            .d       (d),
            .lz      (lz),
            .z       (z)
        );

    end
    else
    begin: POS_EDGE

        mgc_out_reg_pos
        #(
            .rscid   (rscid),
            .width   (width),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        mgc_out_reg_pos_inst
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (ld),
            .d       (d),
            .lz      (lz),
            .z       (z)
        );

    end
    endgenerate

endmodule




//------------------------------------------------------------------

module mgc_out_buf_wait (clk, en, arst, srst, ld, vd, d, vz, lz, z); // Not supported

    parameter integer rscid   = 1;
    parameter integer width   = 8;
    parameter         ph_clk  =  1'b1;
    parameter         ph_en   =  1'b1;
    parameter         ph_arst =  1'b1;
    parameter         ph_srst =  1'b1;

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ld;
    output             vd;
    input  [width-1:0] d;
    output             lz;
    input              vz;
    output [width-1:0] z;

    wire               filled;
    wire               filled_next;
    wire   [width-1:0] abuf;
    wire               lbuf;


    assign filled_next = (filled & (~vz)) | (filled & ld) | (ld & (~vz));

    assign lbuf = ld & ~(filled ^ vz);

    assign vd = vz | ~filled;

    assign lz = ld | filled;

    assign z = (filled) ? abuf : d;

    wire dummy;
    wire dummy_bufreg_lz;

    // Output registers:
    mgc_out_reg
    #(
        .rscid   (rscid),
        .width   (1'b1),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst)
    )
    STATREG
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (filled_next),
        .d       (1'b0),       // input d is unused
        .lz      (filled),
        .z       (dummy)            // output z is unused
    );

    mgc_out_reg
    #(
        .rscid   (rscid),
        .width   (width),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst)
    )
    BUFREG
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (lbuf),
        .d       (d),
        .lz      (dummy_bufreg_lz),
        .z       (abuf)
    );

endmodule

//------------------------------------------------------------------

module mgc_out_fifo_wait (clk, en, arst, srst, ld, vd, d, lz, vz,  z);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer fifo_sz = 8; // fifo depth
    parameter         ph_clk  = 1'b1; // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   = 1'b1; // clock enable polarity
    parameter         ph_arst = 1'b1; // async reset polarity
    parameter         ph_srst = 1'b1; // sync reset polarity
    parameter integer ph_log2 = 3; // log2(fifo_sz)
    parameter integer pwropt  = 0; // pwropt


    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 ld;    // load data
    output                vd;    // fifo full active low
    input     [width-1:0] d;
    output                lz;    // fifo ready to send
    input                 vz;    // dest ready for data
    output    [width-1:0] z;

    wire    [31:0]      size;


      // Output registers:
 mgc_out_fifo_wait_core#(
        .rscid   (rscid),
        .width   (width),
        .sz_width (32),
        .fifo_sz (fifo_sz),
        .ph_clk  (ph_clk),
        .ph_en   (ph_en),
        .ph_arst (ph_arst),
        .ph_srst (ph_srst),
        .ph_log2 (ph_log2),
        .pwropt  (pwropt)
        ) CORE (
        .clk (clk),
        .en (en),
        .arst (arst),
        .srst (srst),
        .ld (ld),
        .vd (vd),
        .d (d),
        .lz (lz),
        .vz (vz),
        .z (z),
        .size (size)
        );

endmodule



module mgc_out_fifo_wait_core (clk, en, arst, srst, ld, vd, d, lz, vz,  z, size);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer sz_width = 8; // size of port for elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter         ph_clk  =  1'b1; // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   =  1'b1; // clock enable polarity
    parameter         ph_arst =  1'b1; // async reset polarity
    parameter         ph_srst =  1'b1; // sync reset polarity
    parameter integer ph_log2 = 3; // log2(fifo_sz)
    parameter integer pwropt  = 0; // pwropt

   localparam integer  fifo_b = width * fifo_sz;

    input                 clk;
    input                 en;
    input                 arst;
    input                 srst;
    input                 ld;    // load data
    output                vd;    // fifo full active low
    input     [width-1:0] d;
    output                lz;    // fifo ready to send
    input                 vz;    // dest ready for data
    output    [width-1:0] z;
    output    [sz_width-1:0]      size;

    reg      [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] stat_pre;
    wire     [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] stat;
    reg      [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff_pre;
    wire     [( (fifo_b > 0) ? fifo_b : 1)-1:0] buff;
    reg      [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] en_l;
    reg      [(((fifo_sz > 0) ? fifo_sz : 1)-1)/8:0] en_l_s;

    reg       [width-1:0] buff_nxt;

    reg                   stat_nxt;
    reg                   stat_before;
    reg                   stat_after;
    reg                   en_l_var;

    integer               i;
    genvar                eni;

    wire [32:0]           size_t;
    reg [31:0]            count;
    reg [31:0]            count_t;
    reg [32:0]            n_elem;
// pragma translate_off
    reg [31:0]            peak;
// pragma translate_on

    wire [( (fifo_sz > 0) ? fifo_sz : 1)-1:0] dummy_statreg_lz;
    wire [( (fifo_b > 0) ? fifo_b : 1)-1:0] dummy_bufreg_lz;

    generate
    if ( fifo_sz > 0 )
    begin: FIFO_REG
      assign vd = vz | ~stat[0];
      assign lz = ld | stat[fifo_sz-1];
      assign size_t = (count - (vz && stat[fifo_sz-1])) + ld;
      assign size = size_t[sz_width-1:0];
      assign z = (stat[fifo_sz-1]) ? buff[fifo_b-1:width*(fifo_sz-1)] : d;

      always @(*)
      begin: FIFOPROC
        n_elem = 33'b0;
        for (i = fifo_sz-1; i >= 0; i = i - 1)
        begin
          if (i != 0)
            stat_before = stat[i-1];
          else
            stat_before = 1'b0;

          if (i != (fifo_sz-1))
            stat_after = stat[i+1];
          else
            stat_after = 1'b1;

          stat_nxt = stat_after &
                    (stat_before | (stat[i] & (~vz)) | (stat[i] & ld) | (ld & (~vz)));

          stat_pre[i] = stat_nxt;
          en_l_var = 1'b1;
          if (!stat_nxt)
            begin
              buff_nxt = {width{1'b0}};
              en_l_var = 1'b0;
            end
          else if (vz && stat_before)
            buff_nxt[0+:width] = buff[width*(i-1)+:width];
          else if (ld && !((vz && stat_before) || ((!vz) && stat[i])))
            buff_nxt = d;
          else
            begin
              if (pwropt == 0)
                buff_nxt[0+:width] = buff[width*i+:width];
              else
                buff_nxt = {width{1'b0}};
              en_l_var = 1'b0;
            end

          if (ph_en != 0)
            en_l[i] = en & en_l_var;
          else
            en_l[i] = en | ~en_l_var;

          buff_pre[width*i+:width] = buff_nxt[0+:width];

          if ((stat_after == 1'b1) && (stat[i] == 1'b0))
            n_elem = ($unsigned(fifo_sz) - 1) - i;
        end

        if (ph_en != 0)
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = 1'b1;
        else
          en_l_s[(((fifo_sz > 0) ? fifo_sz : 1)-1)/8] = 1'b0;

        for (i = fifo_sz-1; i >= 7; i = i - 1)
        begin
          if ((i%'d2) == 0)
          begin
            if (ph_en != 0)
              en_l_s[(i/8)-1] = en & (stat[i]|stat_pre[i-1]);
            else
              en_l_s[(i/8)-1] = en | ~(stat[i]|stat_pre[i-1]);
          end
        end

        if ( stat[fifo_sz-1] == 1'b0 )
          count_t = 32'b0;
        else if ( stat[0] == 1'b1 )
          count_t = { {(32-ph_log2){1'b0}}, fifo_sz};
        else
          count_t = n_elem[31:0];
        count = count_t;
// pragma translate_off
        if ( peak < count )
          peak = count;
// pragma translate_on
      end

      if (pwropt == 0)
      begin: NOCGFIFO
        // Output registers:
        mgc_out_reg
        #(
            .rscid   (rscid),
            .width   (fifo_sz),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        STATREG
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (stat_pre),
            .lz      (dummy_statreg_lz[0]),
            .z       (stat)
        );
        mgc_out_reg
        #(
            .rscid   (rscid),
            .width   (fifo_b),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
        )
        BUFREG
        (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (buff_pre),
            .lz      (dummy_bufreg_lz[0]),
            .z       (buff)
        );
      end
      else
      begin: CGFIFO
        // Output registers:
        if ( pwropt > 1)
        begin: CGSTATFIFO2
          for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
          begin: pwroptGEN1
            mgc_out_reg
            #(
              .rscid   (rscid),
              .width   (1),
              .ph_clk  (ph_clk),
              .ph_en   (ph_en),
              .ph_arst (ph_arst),
              .ph_srst (ph_srst)
            )
            STATREG
            (
              .clk     (clk),
              .en      (en_l_s[eni/8]),
              .arst    (arst),
              .srst    (srst),
              .ld      (1'b1),
              .d       (stat_pre[eni]),
              .lz      (dummy_statreg_lz[eni]),
              .z       (stat[eni])
            );
          end
        end
        else
        begin: CGSTATFIFO
          mgc_out_reg
          #(
            .rscid   (rscid),
            .width   (fifo_sz),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
          )
          STATREG
          (
            .clk     (clk),
            .en      (en),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (stat_pre),
            .lz      (dummy_statreg_lz[0]),
            .z       (stat)
          );
        end
        for (eni = fifo_sz-1; eni >= 0; eni = eni - 1)
        begin: pwroptGEN2
          mgc_out_reg
          #(
            .rscid   (rscid),
            .width   (width),
            .ph_clk  (ph_clk),
            .ph_en   (ph_en),
            .ph_arst (ph_arst),
            .ph_srst (ph_srst)
          )
          BUFREG
          (
            .clk     (clk),
            .en      (en_l[eni]),
            .arst    (arst),
            .srst    (srst),
            .ld      (1'b1),
            .d       (buff_pre[width*eni+:width]),
            .lz      (dummy_bufreg_lz[eni]),
            .z       (buff[width*eni+:width])
          );
        end
      end
    end
    else
    begin: FEED_THRU
      assign vd = vz;
      assign lz = ld;
      assign z = d;
      assign size = ld && !vz;
    end
    endgenerate

endmodule

//------------------------------------------------------------------
//-- PIPE ENTITIES
//------------------------------------------------------------------
/*
 *
 *             _______________________________________________
 * WRITER    |                                               |          READER
 *           |           MGC_PIPE                            |
 *           |           __________________________          |
 *        --<| vdout  --<| vd ---------------  vz<|-----ldin<|---
 *           |           |      FIFO              |          |
 *        ---|>ldout  ---|>ld ---------------- lz |> ---vdin |>--
 *        ---|>dout -----|>d  ---------------- dz |> ----din |>--
 *           |           |________________________|          |
 *           |_______________________________________________|
 */
// two clock pipe
module mgc_pipe (clk, en, arst, srst, ldin, vdin, din, ldout, vdout, dout, size, req_size);

    parameter integer rscid   = 0; // resource ID
    parameter integer width   = 8; // fifo width
    parameter integer sz_width = 8; // width of size of elements in fifo
    parameter integer fifo_sz = 8; // fifo depth
    parameter integer log2_sz = 3; // log2(fifo_sz)
    parameter         ph_clk  = 1'b1;  // clock polarity 1=rising edge, 0=falling edge
    parameter         ph_en   = 1'b1;  // clock enable polarity
    parameter         ph_arst = 1'b1;  // async reset polarity
    parameter         ph_srst = 1'b1;  // sync reset polarity
    parameter integer pwropt  = 0; // pwropt

    input              clk;
    input              en;
    input              arst;
    input              srst;
    input              ldin;
    output             vdin;
    output [width-1:0] din;
    input              ldout;
    output             vdout;
    input  [width-1:0] dout;
    output [sz_width-1:0]      size;
    input              req_size;


    mgc_out_fifo_wait_core
    #(
        .rscid    (rscid),
        .width    (width),
        .sz_width (sz_width),
        .fifo_sz  (fifo_sz),
        .ph_clk   (ph_clk),
        .ph_en    (ph_en),
        .ph_arst  (ph_arst),
        .ph_srst  (ph_srst),
        .ph_log2  (log2_sz),
        .pwropt   (pwropt)
    )
    FIFO
    (
        .clk     (clk),
        .en      (en),
        .arst    (arst),
        .srst    (srst),
        .ld      (ldout),
        .vd      (vdout),
        .d       (dout),
        .lz      (vdin),
        .vz      (ldin),
        .z       (din),
        .size    (size)
    );

endmodule


//------> ./rtl.v 
// ----------------------------------------------------------------------
//  HLS HDL:        Verilog Netlister
//  HLS Version:    2011a.126 Production Release
//  HLS Date:       Wed Aug  8 00:52:07 PDT 2012
// 
//  Generated by:   nn1114@EEWS304-032
//  Generated date: Wed May 13 22:00:42 2015
// ----------------------------------------------------------------------

// 
// ------------------------------------------------------------------
//  Design Unit:    erosion_core_fsm
//  FSM Module
// ------------------------------------------------------------------


module erosion_core_fsm (
  clk, en, arst_n, fsm_output, st_FRAME_tr0
);
  input clk;
  input en;
  input arst_n;
  output [1:0] fsm_output;
  reg [1:0] fsm_output;
  input st_FRAME_tr0;


  // FSM State Type Declaration for erosion_core_fsm_1
  parameter
    st_main = 1'd0,
    st_FRAME = 1'd1,
    state_x = 1'b0;

  reg [0:0] state_var;
  reg [0:0] state_var_NS;


  // Interconnect Declarations for Component Instantiations 
  always @(*)
  begin : erosion_core_fsm_1
    case (state_var)
      st_main : begin
        fsm_output = 2'b1;
        state_var_NS = st_FRAME;
      end
      st_FRAME : begin
        fsm_output = 2'b10;
        if ( st_FRAME_tr0 ) begin
          state_var_NS = st_main;
        end
        else begin
          state_var_NS = st_FRAME;
        end
      end
      default : begin
        fsm_output = 2'b00;
        state_var_NS = st_main;
      end
    endcase
  end

  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      state_var <= st_main;
    end
    else if ( en ) begin
      state_var <= state_var_NS;
    end
  end

endmodule

// ------------------------------------------------------------------
//  Design Unit:    erosion_core
// ------------------------------------------------------------------


module erosion_core (
  clk, en, arst_n, vin_rsc_mgc_in_wire_d, vout_rsc_mgc_out_stdreg_d
);
  input clk;
  input en;
  input arst_n;
  input [149:0] vin_rsc_mgc_in_wire_d;
  output [29:0] vout_rsc_mgc_out_stdreg_d;
  reg [29:0] vout_rsc_mgc_out_stdreg_d;


  // Interconnect Declarations
  wire [1:0] fsm_output;
  wire ACC1_for_nand_tmp;
  wire [2:0] SHIFT_mux_2_tmp;
  wire and_dcpl;
  wire or_dcpl_80;
  wire or_dcpl_83;
  wire or_dcpl_85;
  wire and_dcpl_90;
  wire or_dcpl_93;
  reg apply_lpi_2;
  reg [149:0] regs_operator_din_lpi_2;
  reg exit_SHIFT_lpi_2;
  reg [2:0] ACC1_for_j_1_lpi_2;
  reg [2:0] i_1_lpi_2;
  reg exit_ACC1_lpi_2;
  reg [149:0] regs_regs_0_lpi_2;
  reg [149:0] regs_regs_2_lpi_2;
  reg [149:0] regs_regs_1_lpi_2;
  reg [149:0] regs_regs_3_lpi_2;
  reg [149:0] regs_regs_4_lpi_2;
  reg [18:0] FRAME_p_1_sva;
  reg exit_ACC1_1_sva;
  reg exit_ACC1_for_lpi_2_dfm_1;
  reg [149:0] regs_regs_0_lpi_2_dfm_1;
  reg [149:0] regs_regs_1_lpi_2_dfm_1;
  reg [149:0] regs_regs_2_lpi_2_dfm_1;
  reg [149:0] regs_regs_3_lpi_2_dfm_1;
  reg [149:0] regs_regs_4_lpi_2_dfm_1;
  reg apply_lpi_2_dfm_2;
  reg [2:0] i_1_lpi_2_dfm_2;
  reg [2:0] ACC1_for_j_1_lpi_2_dfm_4;
  reg exit_ACC1_lpi_2_dfm_3;
  reg exit_SHIFT_lpi_2_dfm_1;
  reg FRAME_stage_0;
  reg [2:0] SHIFT_i_1_lpi_5;
  wire and_89_cse;
  wire and_88_cse;
  wire exit_SHIFT_lpi_2_dfm_2;
  wire [2:0] SHIFT_acc_1_psp;
  wire [3:0] nl_SHIFT_acc_1_psp;
  wire or_dcpl_113;
  wire and_dcpl_136;
  wire or_dcpl_115;
  wire or_dcpl_116;
  wire SHIFT_and_8_cse;
  wire nor_8_cse;
  wire SHIFT_and_cse;
  wire [2:0] ACC1_for_acc_itm;
  wire [3:0] nl_ACC1_for_acc_itm;
  wire [2:0] ACC1_acc_itm;
  wire [3:0] nl_ACC1_acc_itm;
  wire [2:0] i_1_lpi_2_dfm_2_mx1w0;
  wire [2:0] ACC1_for_j_1_lpi_2_dfm_4_mx1w0;
  wire exit_ACC1_for_lpi_2_dfm_1_mx2;
  wire [149:0] regs_operator_din_lpi_2_mx0;
  wire [18:0] FRAME_p_1_sva_1;
  wire [19:0] nl_FRAME_p_1_sva_1;
  wire apply_lpi_2_dfm_1;
  wire exit_ACC1_lpi_2_dfm_1_mx0;
  wire [2:0] i_1_sva;
  wire [3:0] nl_i_1_sva;
  wire [2:0] ACC1_for_j_1_sva;
  wire [3:0] nl_ACC1_for_j_1_sva;
  wire apply_lpi_2_dfm;
  wire [1:0] ACC1_for_slc_1_svs_sg14;
  wire [1:0] ACC1_for_slc_1_svs_sg13;
  wire [1:0] ACC1_for_slc_1_svs_sg12;
  wire [1:0] ACC1_for_slc_1_svs_sg11;
  wire [1:0] ACC1_for_slc_1_svs_sg10;
  wire [1:0] ACC1_for_slc_1_svs_sg9;
  wire [1:0] ACC1_for_slc_1_svs_sg8;
  wire [1:0] ACC1_for_slc_1_svs_sg7;
  wire [1:0] ACC1_for_slc_1_svs_sg6;
  wire [1:0] ACC1_for_slc_1_svs_sg5;
  wire [1:0] ACC1_for_slc_1_svs_sg4;
  wire [1:0] ACC1_for_slc_1_svs_sg3;
  wire [1:0] ACC1_for_slc_1_svs_sg2;
  wire [1:0] ACC1_for_slc_1_svs_sg1;
  wire [1:0] ACC1_for_slc_1_svs_1;
  wire [8:0] ACC1_for_if_acc_ssc;
  wire [9:0] nl_ACC1_for_if_acc_ssc;
  wire [2:0] SHIFT_i_1_lpi_2_dfm_2_mx0;
  wire [149:0] SHIFT_if_else_else_else_slc_regs_regs_ctmp_sva;
  wire and_151_cse;
  wire and_152_cse;

  wire[2:0] mux_25_nl;
  wire[2:0] mux_26_nl;
  wire[0:0] mux_nl;

  // Interconnect Declarations for Component Instantiations 
  wire [0:0] nl_erosion_core_fsm_inst_st_FRAME_tr0;
  assign nl_erosion_core_fsm_inst_st_FRAME_tr0 = ~ FRAME_stage_0;
  erosion_core_fsm erosion_core_fsm_inst (
      .clk(clk),
      .en(en),
      .arst_n(arst_n),
      .fsm_output(fsm_output),
      .st_FRAME_tr0(nl_erosion_core_fsm_inst_st_FRAME_tr0)
    );
  assign and_151_cse = (~ FRAME_stage_0) & (fsm_output[1]);
  assign and_152_cse = FRAME_stage_0 & (fsm_output[1]);
  assign mux_25_nl = MUX_v_3_2_2({i_1_sva , i_1_lpi_2}, or_dcpl_113);
  assign i_1_lpi_2_dfm_2_mx1w0 = ~((~((mux_25_nl) | (signext_3_1(~(SHIFT_and_8_cse
      | or_dcpl_113 | and_dcpl_136))))) | ({{2{and_dcpl_136}}, and_dcpl_136}));
  assign mux_26_nl = MUX_v_3_2_2({ACC1_for_j_1_sva , ACC1_for_j_1_lpi_2}, or_dcpl_115);
  assign ACC1_for_j_1_lpi_2_dfm_4_mx1w0 = ~((~((mux_26_nl) | (signext_3_1(~((SHIFT_and_8_cse
      & (~ ACC1_for_nand_tmp) & (~ (ACC1_acc_itm[2]))) | SHIFT_and_cse | or_dcpl_115
      | or_dcpl_116))))) | ({{2{or_dcpl_116}}, or_dcpl_116}));
  assign nl_ACC1_for_acc_itm = ACC1_for_j_1_sva + 3'b11;
  assign ACC1_for_acc_itm = nl_ACC1_for_acc_itm[2:0];
  assign mux_nl = MUX_s_1_2_2({(~ (ACC1_for_acc_itm[2])) , exit_ACC1_for_lpi_2_dfm_1},
      or_dcpl_80);
  assign exit_ACC1_for_lpi_2_dfm_1_mx2 = (mux_nl) | (exit_SHIFT_lpi_2_dfm_2 & ACC1_for_nand_tmp);
  assign regs_operator_din_lpi_2_mx0 = MUX_v_150_2_2({regs_operator_din_lpi_2 , vin_rsc_mgc_in_wire_d},
      exit_ACC1_1_sva);
  assign nl_FRAME_p_1_sva_1 = FRAME_p_1_sva + 19'b1;
  assign FRAME_p_1_sva_1 = nl_FRAME_p_1_sva_1[18:0];
  assign apply_lpi_2_dfm_1 = apply_lpi_2_dfm & (~ ACC1_for_nand_tmp);
  assign exit_ACC1_lpi_2_dfm_1_mx0 = MUX_s_1_2_2({(~ (ACC1_acc_itm[2])) , exit_ACC1_lpi_2},
      and_dcpl);
  assign nl_ACC1_acc_itm = i_1_sva + 3'b11;
  assign ACC1_acc_itm = nl_ACC1_acc_itm[2:0];
  assign nl_i_1_sva = i_1_lpi_2 + 3'b1;
  assign i_1_sva = nl_i_1_sva[2:0];
  assign nl_ACC1_for_j_1_sva = ACC1_for_j_1_lpi_2 + 3'b1;
  assign ACC1_for_j_1_sva = nl_ACC1_for_j_1_sva[2:0];
  assign ACC1_for_nand_tmp = ~((ACC1_for_slc_1_svs_sg14[1]) & (ACC1_for_slc_1_svs_sg14[0])
      & (ACC1_for_slc_1_svs_sg13[1]) & (ACC1_for_slc_1_svs_sg13[0]) & (ACC1_for_slc_1_svs_sg12[1])
      & (ACC1_for_slc_1_svs_sg12[0]) & (ACC1_for_slc_1_svs_sg11[1]) & (ACC1_for_slc_1_svs_sg11[0])
      & (ACC1_for_slc_1_svs_sg10[1]) & (ACC1_for_slc_1_svs_sg10[0]) & (ACC1_for_slc_1_svs_sg9[1])
      & (ACC1_for_slc_1_svs_sg9[0]) & (ACC1_for_slc_1_svs_sg8[1]) & (ACC1_for_slc_1_svs_sg8[0])
      & (ACC1_for_slc_1_svs_sg7[1]) & (ACC1_for_slc_1_svs_sg7[0]) & (ACC1_for_slc_1_svs_sg6[1])
      & (ACC1_for_slc_1_svs_sg6[0]) & (ACC1_for_slc_1_svs_sg5[1]) & (ACC1_for_slc_1_svs_sg5[0])
      & (ACC1_for_slc_1_svs_sg4[1]) & (ACC1_for_slc_1_svs_sg4[0]) & (ACC1_for_slc_1_svs_sg3[1])
      & (ACC1_for_slc_1_svs_sg3[0]) & (ACC1_for_slc_1_svs_sg2[1]) & (ACC1_for_slc_1_svs_sg2[0])
      & (ACC1_for_slc_1_svs_sg1[1]) & (ACC1_for_slc_1_svs_sg1[0]) & (ACC1_for_slc_1_svs_1[1])
      & (ACC1_for_slc_1_svs_1[0]));
  assign apply_lpi_2_dfm = apply_lpi_2 | exit_ACC1_1_sva;
  assign ACC1_for_slc_1_svs_sg14 = MUX_v_2_512_2({(regs_regs_0_lpi_2[29:28]) , (regs_regs_0_lpi_2[31:30])
      , (regs_regs_0_lpi_2[33:32]) , (regs_regs_0_lpi_2[35:34]) , (regs_regs_0_lpi_2[37:36])
      , (regs_regs_0_lpi_2[39:38]) , (regs_regs_0_lpi_2[41:40]) , (regs_regs_0_lpi_2[43:42])
      , (regs_regs_0_lpi_2[45:44]) , (regs_regs_0_lpi_2[47:46]) , (regs_regs_0_lpi_2[49:48])
      , (regs_regs_0_lpi_2[51:50]) , (regs_regs_0_lpi_2[53:52]) , (regs_regs_0_lpi_2[55:54])
      , (regs_regs_0_lpi_2[57:56]) , (regs_regs_0_lpi_2[59:58]) , (regs_regs_0_lpi_2[61:60])
      , (regs_regs_0_lpi_2[63:62]) , (regs_regs_0_lpi_2[65:64]) , (regs_regs_0_lpi_2[67:66])
      , (regs_regs_0_lpi_2[69:68]) , (regs_regs_0_lpi_2[71:70]) , (regs_regs_0_lpi_2[73:72])
      , (regs_regs_0_lpi_2[75:74]) , (regs_regs_0_lpi_2[77:76]) , (regs_regs_0_lpi_2[79:78])
      , (regs_regs_0_lpi_2[81:80]) , (regs_regs_0_lpi_2[83:82]) , (regs_regs_0_lpi_2[85:84])
      , (regs_regs_0_lpi_2[87:86]) , (regs_regs_0_lpi_2[89:88]) , (regs_regs_0_lpi_2[91:90])
      , (regs_regs_0_lpi_2[93:92]) , (regs_regs_0_lpi_2[95:94]) , (regs_regs_0_lpi_2[97:96])
      , (regs_regs_0_lpi_2[99:98]) , (regs_regs_0_lpi_2[101:100]) , (regs_regs_0_lpi_2[103:102])
      , (regs_regs_0_lpi_2[105:104]) , (regs_regs_0_lpi_2[107:106]) , (regs_regs_0_lpi_2[109:108])
      , (regs_regs_0_lpi_2[111:110]) , (regs_regs_0_lpi_2[113:112]) , (regs_regs_0_lpi_2[115:114])
      , (regs_regs_0_lpi_2[117:116]) , (regs_regs_0_lpi_2[119:118]) , (regs_regs_0_lpi_2[121:120])
      , (regs_regs_0_lpi_2[123:122]) , (regs_regs_0_lpi_2[125:124]) , (regs_regs_0_lpi_2[127:126])
      , (regs_regs_0_lpi_2[129:128]) , (regs_regs_0_lpi_2[131:130]) , (regs_regs_0_lpi_2[133:132])
      , (regs_regs_0_lpi_2[135:134]) , (regs_regs_0_lpi_2[137:136]) , (regs_regs_0_lpi_2[139:138])
      , (regs_regs_0_lpi_2[141:140]) , (regs_regs_0_lpi_2[143:142]) , (regs_regs_0_lpi_2[145:144])
      , (regs_regs_0_lpi_2[147:146]) , (regs_regs_0_lpi_2[149:148]) , (regs_regs_1_lpi_2[1:0])
      , (regs_regs_1_lpi_2[3:2]) , (regs_regs_1_lpi_2[5:4]) , (regs_regs_1_lpi_2[7:6])
      , (regs_regs_1_lpi_2[9:8]) , (regs_regs_1_lpi_2[11:10]) , (regs_regs_1_lpi_2[13:12])
      , (regs_regs_1_lpi_2[15:14]) , (regs_regs_1_lpi_2[17:16]) , (regs_regs_1_lpi_2[19:18])
      , (regs_regs_1_lpi_2[21:20]) , (regs_regs_1_lpi_2[23:22]) , (regs_regs_1_lpi_2[25:24])
      , (regs_regs_1_lpi_2[27:26]) , (regs_regs_1_lpi_2[29:28]) , (regs_regs_1_lpi_2[31:30])
      , (regs_regs_1_lpi_2[33:32]) , (regs_regs_1_lpi_2[35:34]) , (regs_regs_1_lpi_2[37:36])
      , (regs_regs_1_lpi_2[39:38]) , (regs_regs_1_lpi_2[41:40]) , (regs_regs_1_lpi_2[43:42])
      , (regs_regs_1_lpi_2[45:44]) , (regs_regs_1_lpi_2[47:46]) , (regs_regs_1_lpi_2[49:48])
      , (regs_regs_1_lpi_2[51:50]) , (regs_regs_1_lpi_2[53:52]) , (regs_regs_1_lpi_2[55:54])
      , (regs_regs_1_lpi_2[57:56]) , (regs_regs_1_lpi_2[59:58]) , (regs_regs_1_lpi_2[61:60])
      , (regs_regs_1_lpi_2[63:62]) , (regs_regs_1_lpi_2[65:64]) , (regs_regs_1_lpi_2[67:66])
      , (regs_regs_1_lpi_2[69:68]) , (regs_regs_1_lpi_2[71:70]) , (regs_regs_1_lpi_2[73:72])
      , (regs_regs_1_lpi_2[75:74]) , (regs_regs_1_lpi_2[77:76]) , (regs_regs_1_lpi_2[79:78])
      , (regs_regs_1_lpi_2[81:80]) , (regs_regs_1_lpi_2[83:82]) , (regs_regs_1_lpi_2[85:84])
      , (regs_regs_1_lpi_2[87:86]) , (regs_regs_1_lpi_2[89:88]) , (regs_regs_1_lpi_2[91:90])
      , (regs_regs_1_lpi_2[93:92]) , (regs_regs_1_lpi_2[95:94]) , (regs_regs_1_lpi_2[97:96])
      , (regs_regs_1_lpi_2[99:98]) , (regs_regs_1_lpi_2[101:100]) , (regs_regs_1_lpi_2[103:102])
      , (regs_regs_1_lpi_2[105:104]) , (regs_regs_1_lpi_2[107:106]) , (regs_regs_1_lpi_2[109:108])
      , (regs_regs_1_lpi_2[111:110]) , (regs_regs_1_lpi_2[113:112]) , (regs_regs_1_lpi_2[115:114])
      , (regs_regs_1_lpi_2[117:116]) , (regs_regs_1_lpi_2[119:118]) , (regs_regs_1_lpi_2[121:120])
      , (regs_regs_1_lpi_2[123:122]) , (regs_regs_1_lpi_2[125:124]) , (regs_regs_1_lpi_2[127:126])
      , (regs_regs_1_lpi_2[129:128]) , (regs_regs_1_lpi_2[131:130]) , (regs_regs_1_lpi_2[133:132])
      , (regs_regs_1_lpi_2[135:134]) , (regs_regs_1_lpi_2[137:136]) , (regs_regs_1_lpi_2[139:138])
      , (regs_regs_1_lpi_2[141:140]) , (regs_regs_1_lpi_2[143:142]) , (regs_regs_1_lpi_2[145:144])
      , (regs_regs_1_lpi_2[147:146]) , (regs_regs_1_lpi_2[149:148]) , (regs_regs_2_lpi_2[1:0])
      , (regs_regs_2_lpi_2[3:2]) , (regs_regs_2_lpi_2[5:4]) , (regs_regs_2_lpi_2[7:6])
      , (regs_regs_2_lpi_2[9:8]) , (regs_regs_2_lpi_2[11:10]) , (regs_regs_2_lpi_2[13:12])
      , (regs_regs_2_lpi_2[15:14]) , (regs_regs_2_lpi_2[17:16]) , (regs_regs_2_lpi_2[19:18])
      , (regs_regs_2_lpi_2[21:20]) , (regs_regs_2_lpi_2[23:22]) , (regs_regs_2_lpi_2[25:24])
      , (regs_regs_2_lpi_2[27:26]) , (regs_regs_2_lpi_2[29:28]) , (regs_regs_2_lpi_2[31:30])
      , (regs_regs_2_lpi_2[33:32]) , (regs_regs_2_lpi_2[35:34]) , (regs_regs_2_lpi_2[37:36])
      , (regs_regs_2_lpi_2[39:38]) , (regs_regs_2_lpi_2[41:40]) , (regs_regs_2_lpi_2[43:42])
      , (regs_regs_2_lpi_2[45:44]) , (regs_regs_2_lpi_2[47:46]) , (regs_regs_2_lpi_2[49:48])
      , (regs_regs_2_lpi_2[51:50]) , (regs_regs_2_lpi_2[53:52]) , (regs_regs_2_lpi_2[55:54])
      , (regs_regs_2_lpi_2[57:56]) , (regs_regs_2_lpi_2[59:58]) , (regs_regs_2_lpi_2[61:60])
      , (regs_regs_2_lpi_2[63:62]) , (regs_regs_2_lpi_2[65:64]) , (regs_regs_2_lpi_2[67:66])
      , (regs_regs_2_lpi_2[69:68]) , (regs_regs_2_lpi_2[71:70]) , (regs_regs_2_lpi_2[73:72])
      , (regs_regs_2_lpi_2[75:74]) , (regs_regs_2_lpi_2[77:76]) , (regs_regs_2_lpi_2[79:78])
      , (regs_regs_2_lpi_2[81:80]) , (regs_regs_2_lpi_2[83:82]) , (regs_regs_2_lpi_2[85:84])
      , (regs_regs_2_lpi_2[87:86]) , (regs_regs_2_lpi_2[89:88]) , (regs_regs_2_lpi_2[91:90])
      , (regs_regs_2_lpi_2[93:92]) , (regs_regs_2_lpi_2[95:94]) , (regs_regs_2_lpi_2[97:96])
      , (regs_regs_2_lpi_2[99:98]) , (regs_regs_2_lpi_2[101:100]) , (regs_regs_2_lpi_2[103:102])
      , (regs_regs_2_lpi_2[105:104]) , (regs_regs_2_lpi_2[107:106]) , (regs_regs_2_lpi_2[109:108])
      , (regs_regs_2_lpi_2[111:110]) , (regs_regs_2_lpi_2[113:112]) , (regs_regs_2_lpi_2[115:114])
      , (regs_regs_2_lpi_2[117:116]) , (regs_regs_2_lpi_2[119:118]) , (regs_regs_2_lpi_2[121:120])
      , (regs_regs_2_lpi_2[123:122]) , (regs_regs_2_lpi_2[125:124]) , (regs_regs_2_lpi_2[127:126])
      , (regs_regs_2_lpi_2[129:128]) , (regs_regs_2_lpi_2[131:130]) , (regs_regs_2_lpi_2[133:132])
      , (regs_regs_2_lpi_2[135:134]) , (regs_regs_2_lpi_2[137:136]) , (regs_regs_2_lpi_2[139:138])
      , (regs_regs_2_lpi_2[141:140]) , (regs_regs_2_lpi_2[143:142]) , (regs_regs_2_lpi_2[145:144])
      , (regs_regs_2_lpi_2[147:146]) , (regs_regs_2_lpi_2[149:148]) , (regs_regs_3_lpi_2[1:0])
      , (regs_regs_3_lpi_2[3:2]) , (regs_regs_3_lpi_2[5:4]) , (regs_regs_3_lpi_2[7:6])
      , (regs_regs_3_lpi_2[9:8]) , (regs_regs_3_lpi_2[11:10]) , (regs_regs_3_lpi_2[13:12])
      , (regs_regs_3_lpi_2[15:14]) , (regs_regs_3_lpi_2[17:16]) , (regs_regs_3_lpi_2[19:18])
      , (regs_regs_3_lpi_2[21:20]) , (regs_regs_3_lpi_2[23:22]) , (regs_regs_3_lpi_2[25:24])
      , (regs_regs_3_lpi_2[27:26]) , (regs_regs_3_lpi_2[29:28]) , (regs_regs_3_lpi_2[31:30])
      , (regs_regs_3_lpi_2[33:32]) , (regs_regs_3_lpi_2[35:34]) , (regs_regs_3_lpi_2[37:36])
      , (regs_regs_3_lpi_2[39:38]) , (regs_regs_3_lpi_2[41:40]) , (regs_regs_3_lpi_2[43:42])
      , (regs_regs_3_lpi_2[45:44]) , (regs_regs_3_lpi_2[47:46]) , (regs_regs_3_lpi_2[49:48])
      , (regs_regs_3_lpi_2[51:50]) , (regs_regs_3_lpi_2[53:52]) , (regs_regs_3_lpi_2[55:54])
      , (regs_regs_3_lpi_2[57:56]) , (regs_regs_3_lpi_2[59:58]) , (regs_regs_3_lpi_2[61:60])
      , (regs_regs_3_lpi_2[63:62]) , (regs_regs_3_lpi_2[65:64]) , (regs_regs_3_lpi_2[67:66])
      , (regs_regs_3_lpi_2[69:68]) , (regs_regs_3_lpi_2[71:70]) , (regs_regs_3_lpi_2[73:72])
      , (regs_regs_3_lpi_2[75:74]) , (regs_regs_3_lpi_2[77:76]) , (regs_regs_3_lpi_2[79:78])
      , (regs_regs_3_lpi_2[81:80]) , (regs_regs_3_lpi_2[83:82]) , (regs_regs_3_lpi_2[85:84])
      , (regs_regs_3_lpi_2[87:86]) , (regs_regs_3_lpi_2[89:88]) , (regs_regs_3_lpi_2[91:90])
      , (regs_regs_3_lpi_2[93:92]) , (regs_regs_3_lpi_2[95:94]) , (regs_regs_3_lpi_2[97:96])
      , (regs_regs_3_lpi_2[99:98]) , (regs_regs_3_lpi_2[101:100]) , (regs_regs_3_lpi_2[103:102])
      , (regs_regs_3_lpi_2[105:104]) , (regs_regs_3_lpi_2[107:106]) , (regs_regs_3_lpi_2[109:108])
      , (regs_regs_3_lpi_2[111:110]) , (regs_regs_3_lpi_2[113:112]) , (regs_regs_3_lpi_2[115:114])
      , (regs_regs_3_lpi_2[117:116]) , (regs_regs_3_lpi_2[119:118]) , (regs_regs_3_lpi_2[121:120])
      , (regs_regs_3_lpi_2[123:122]) , (regs_regs_3_lpi_2[125:124]) , (regs_regs_3_lpi_2[127:126])
      , (regs_regs_3_lpi_2[129:128]) , (regs_regs_3_lpi_2[131:130]) , (regs_regs_3_lpi_2[133:132])
      , (regs_regs_3_lpi_2[135:134]) , (regs_regs_3_lpi_2[137:136]) , (regs_regs_3_lpi_2[139:138])
      , (regs_regs_3_lpi_2[141:140]) , (regs_regs_3_lpi_2[143:142]) , (regs_regs_3_lpi_2[145:144])
      , (regs_regs_3_lpi_2[147:146]) , (regs_regs_3_lpi_2[149:148]) , (regs_regs_4_lpi_2[1:0])
      , (regs_regs_4_lpi_2[3:2]) , (regs_regs_4_lpi_2[5:4]) , (regs_regs_4_lpi_2[7:6])
      , (regs_regs_4_lpi_2[9:8]) , (regs_regs_4_lpi_2[11:10]) , (regs_regs_4_lpi_2[13:12])
      , (regs_regs_4_lpi_2[15:14]) , (regs_regs_4_lpi_2[17:16]) , (regs_regs_4_lpi_2[19:18])
      , (regs_regs_4_lpi_2[21:20]) , (regs_regs_4_lpi_2[23:22]) , (regs_regs_4_lpi_2[25:24])
      , (regs_regs_4_lpi_2[27:26]) , (regs_regs_4_lpi_2[29:28]) , (regs_regs_4_lpi_2[31:30])
      , (regs_regs_4_lpi_2[33:32]) , (regs_regs_4_lpi_2[35:34]) , (regs_regs_4_lpi_2[37:36])
      , (regs_regs_4_lpi_2[39:38]) , (regs_regs_4_lpi_2[41:40]) , (regs_regs_4_lpi_2[43:42])
      , (regs_regs_4_lpi_2[45:44]) , (regs_regs_4_lpi_2[47:46]) , (regs_regs_4_lpi_2[49:48])
      , (regs_regs_4_lpi_2[51:50]) , (regs_regs_4_lpi_2[53:52]) , (regs_regs_4_lpi_2[55:54])
      , (regs_regs_4_lpi_2[57:56]) , (regs_regs_4_lpi_2[59:58]) , (regs_regs_4_lpi_2[61:60])
      , (regs_regs_4_lpi_2[63:62]) , (regs_regs_4_lpi_2[65:64]) , (regs_regs_4_lpi_2[67:66])
      , (regs_regs_4_lpi_2[69:68]) , (regs_regs_4_lpi_2[71:70]) , (regs_regs_4_lpi_2[73:72])
      , (regs_regs_4_lpi_2[75:74]) , (regs_regs_4_lpi_2[77:76]) , (regs_regs_4_lpi_2[79:78])
      , (regs_regs_4_lpi_2[81:80]) , (regs_regs_4_lpi_2[83:82]) , (regs_regs_4_lpi_2[85:84])
      , (regs_regs_4_lpi_2[87:86]) , (regs_regs_4_lpi_2[89:88]) , (regs_regs_4_lpi_2[91:90])
      , (regs_regs_4_lpi_2[93:92]) , (regs_regs_4_lpi_2[95:94]) , (regs_regs_4_lpi_2[97:96])
      , (regs_regs_4_lpi_2[99:98]) , (regs_regs_4_lpi_2[101:100]) , (regs_regs_4_lpi_2[103:102])
      , (regs_regs_4_lpi_2[105:104]) , (regs_regs_4_lpi_2[107:106]) , (regs_regs_4_lpi_2[109:108])
      , (regs_regs_4_lpi_2[111:110]) , (regs_regs_4_lpi_2[113:112]) , (regs_regs_4_lpi_2[115:114])
      , (regs_regs_4_lpi_2[117:116]) , (regs_regs_4_lpi_2[119:118]) , (regs_regs_4_lpi_2[121:120])
      , (regs_regs_4_lpi_2[123:122]) , (regs_regs_4_lpi_2[125:124]) , (regs_regs_4_lpi_2[127:126])
      , (regs_regs_4_lpi_2[129:128]) , (regs_regs_4_lpi_2[131:130]) , (regs_regs_4_lpi_2[133:132])
      , (regs_regs_4_lpi_2[135:134]) , (regs_regs_4_lpi_2[137:136]) , (regs_regs_4_lpi_2[139:138])
      , (regs_regs_4_lpi_2[141:140]) , (regs_regs_4_lpi_2[143:142]) , (regs_regs_4_lpi_2[145:144])
      , (regs_regs_4_lpi_2[147:146]) , (regs_regs_4_lpi_2[149:148]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg13 = MUX_v_2_512_2({(regs_regs_0_lpi_2[27:26]) , (regs_regs_0_lpi_2[29:28])
      , (regs_regs_0_lpi_2[31:30]) , (regs_regs_0_lpi_2[33:32]) , (regs_regs_0_lpi_2[35:34])
      , (regs_regs_0_lpi_2[37:36]) , (regs_regs_0_lpi_2[39:38]) , (regs_regs_0_lpi_2[41:40])
      , (regs_regs_0_lpi_2[43:42]) , (regs_regs_0_lpi_2[45:44]) , (regs_regs_0_lpi_2[47:46])
      , (regs_regs_0_lpi_2[49:48]) , (regs_regs_0_lpi_2[51:50]) , (regs_regs_0_lpi_2[53:52])
      , (regs_regs_0_lpi_2[55:54]) , (regs_regs_0_lpi_2[57:56]) , (regs_regs_0_lpi_2[59:58])
      , (regs_regs_0_lpi_2[61:60]) , (regs_regs_0_lpi_2[63:62]) , (regs_regs_0_lpi_2[65:64])
      , (regs_regs_0_lpi_2[67:66]) , (regs_regs_0_lpi_2[69:68]) , (regs_regs_0_lpi_2[71:70])
      , (regs_regs_0_lpi_2[73:72]) , (regs_regs_0_lpi_2[75:74]) , (regs_regs_0_lpi_2[77:76])
      , (regs_regs_0_lpi_2[79:78]) , (regs_regs_0_lpi_2[81:80]) , (regs_regs_0_lpi_2[83:82])
      , (regs_regs_0_lpi_2[85:84]) , (regs_regs_0_lpi_2[87:86]) , (regs_regs_0_lpi_2[89:88])
      , (regs_regs_0_lpi_2[91:90]) , (regs_regs_0_lpi_2[93:92]) , (regs_regs_0_lpi_2[95:94])
      , (regs_regs_0_lpi_2[97:96]) , (regs_regs_0_lpi_2[99:98]) , (regs_regs_0_lpi_2[101:100])
      , (regs_regs_0_lpi_2[103:102]) , (regs_regs_0_lpi_2[105:104]) , (regs_regs_0_lpi_2[107:106])
      , (regs_regs_0_lpi_2[109:108]) , (regs_regs_0_lpi_2[111:110]) , (regs_regs_0_lpi_2[113:112])
      , (regs_regs_0_lpi_2[115:114]) , (regs_regs_0_lpi_2[117:116]) , (regs_regs_0_lpi_2[119:118])
      , (regs_regs_0_lpi_2[121:120]) , (regs_regs_0_lpi_2[123:122]) , (regs_regs_0_lpi_2[125:124])
      , (regs_regs_0_lpi_2[127:126]) , (regs_regs_0_lpi_2[129:128]) , (regs_regs_0_lpi_2[131:130])
      , (regs_regs_0_lpi_2[133:132]) , (regs_regs_0_lpi_2[135:134]) , (regs_regs_0_lpi_2[137:136])
      , (regs_regs_0_lpi_2[139:138]) , (regs_regs_0_lpi_2[141:140]) , (regs_regs_0_lpi_2[143:142])
      , (regs_regs_0_lpi_2[145:144]) , (regs_regs_0_lpi_2[147:146]) , (regs_regs_0_lpi_2[149:148])
      , (regs_regs_1_lpi_2[1:0]) , (regs_regs_1_lpi_2[3:2]) , (regs_regs_1_lpi_2[5:4])
      , (regs_regs_1_lpi_2[7:6]) , (regs_regs_1_lpi_2[9:8]) , (regs_regs_1_lpi_2[11:10])
      , (regs_regs_1_lpi_2[13:12]) , (regs_regs_1_lpi_2[15:14]) , (regs_regs_1_lpi_2[17:16])
      , (regs_regs_1_lpi_2[19:18]) , (regs_regs_1_lpi_2[21:20]) , (regs_regs_1_lpi_2[23:22])
      , (regs_regs_1_lpi_2[25:24]) , (regs_regs_1_lpi_2[27:26]) , (regs_regs_1_lpi_2[29:28])
      , (regs_regs_1_lpi_2[31:30]) , (regs_regs_1_lpi_2[33:32]) , (regs_regs_1_lpi_2[35:34])
      , (regs_regs_1_lpi_2[37:36]) , (regs_regs_1_lpi_2[39:38]) , (regs_regs_1_lpi_2[41:40])
      , (regs_regs_1_lpi_2[43:42]) , (regs_regs_1_lpi_2[45:44]) , (regs_regs_1_lpi_2[47:46])
      , (regs_regs_1_lpi_2[49:48]) , (regs_regs_1_lpi_2[51:50]) , (regs_regs_1_lpi_2[53:52])
      , (regs_regs_1_lpi_2[55:54]) , (regs_regs_1_lpi_2[57:56]) , (regs_regs_1_lpi_2[59:58])
      , (regs_regs_1_lpi_2[61:60]) , (regs_regs_1_lpi_2[63:62]) , (regs_regs_1_lpi_2[65:64])
      , (regs_regs_1_lpi_2[67:66]) , (regs_regs_1_lpi_2[69:68]) , (regs_regs_1_lpi_2[71:70])
      , (regs_regs_1_lpi_2[73:72]) , (regs_regs_1_lpi_2[75:74]) , (regs_regs_1_lpi_2[77:76])
      , (regs_regs_1_lpi_2[79:78]) , (regs_regs_1_lpi_2[81:80]) , (regs_regs_1_lpi_2[83:82])
      , (regs_regs_1_lpi_2[85:84]) , (regs_regs_1_lpi_2[87:86]) , (regs_regs_1_lpi_2[89:88])
      , (regs_regs_1_lpi_2[91:90]) , (regs_regs_1_lpi_2[93:92]) , (regs_regs_1_lpi_2[95:94])
      , (regs_regs_1_lpi_2[97:96]) , (regs_regs_1_lpi_2[99:98]) , (regs_regs_1_lpi_2[101:100])
      , (regs_regs_1_lpi_2[103:102]) , (regs_regs_1_lpi_2[105:104]) , (regs_regs_1_lpi_2[107:106])
      , (regs_regs_1_lpi_2[109:108]) , (regs_regs_1_lpi_2[111:110]) , (regs_regs_1_lpi_2[113:112])
      , (regs_regs_1_lpi_2[115:114]) , (regs_regs_1_lpi_2[117:116]) , (regs_regs_1_lpi_2[119:118])
      , (regs_regs_1_lpi_2[121:120]) , (regs_regs_1_lpi_2[123:122]) , (regs_regs_1_lpi_2[125:124])
      , (regs_regs_1_lpi_2[127:126]) , (regs_regs_1_lpi_2[129:128]) , (regs_regs_1_lpi_2[131:130])
      , (regs_regs_1_lpi_2[133:132]) , (regs_regs_1_lpi_2[135:134]) , (regs_regs_1_lpi_2[137:136])
      , (regs_regs_1_lpi_2[139:138]) , (regs_regs_1_lpi_2[141:140]) , (regs_regs_1_lpi_2[143:142])
      , (regs_regs_1_lpi_2[145:144]) , (regs_regs_1_lpi_2[147:146]) , (regs_regs_1_lpi_2[149:148])
      , (regs_regs_2_lpi_2[1:0]) , (regs_regs_2_lpi_2[3:2]) , (regs_regs_2_lpi_2[5:4])
      , (regs_regs_2_lpi_2[7:6]) , (regs_regs_2_lpi_2[9:8]) , (regs_regs_2_lpi_2[11:10])
      , (regs_regs_2_lpi_2[13:12]) , (regs_regs_2_lpi_2[15:14]) , (regs_regs_2_lpi_2[17:16])
      , (regs_regs_2_lpi_2[19:18]) , (regs_regs_2_lpi_2[21:20]) , (regs_regs_2_lpi_2[23:22])
      , (regs_regs_2_lpi_2[25:24]) , (regs_regs_2_lpi_2[27:26]) , (regs_regs_2_lpi_2[29:28])
      , (regs_regs_2_lpi_2[31:30]) , (regs_regs_2_lpi_2[33:32]) , (regs_regs_2_lpi_2[35:34])
      , (regs_regs_2_lpi_2[37:36]) , (regs_regs_2_lpi_2[39:38]) , (regs_regs_2_lpi_2[41:40])
      , (regs_regs_2_lpi_2[43:42]) , (regs_regs_2_lpi_2[45:44]) , (regs_regs_2_lpi_2[47:46])
      , (regs_regs_2_lpi_2[49:48]) , (regs_regs_2_lpi_2[51:50]) , (regs_regs_2_lpi_2[53:52])
      , (regs_regs_2_lpi_2[55:54]) , (regs_regs_2_lpi_2[57:56]) , (regs_regs_2_lpi_2[59:58])
      , (regs_regs_2_lpi_2[61:60]) , (regs_regs_2_lpi_2[63:62]) , (regs_regs_2_lpi_2[65:64])
      , (regs_regs_2_lpi_2[67:66]) , (regs_regs_2_lpi_2[69:68]) , (regs_regs_2_lpi_2[71:70])
      , (regs_regs_2_lpi_2[73:72]) , (regs_regs_2_lpi_2[75:74]) , (regs_regs_2_lpi_2[77:76])
      , (regs_regs_2_lpi_2[79:78]) , (regs_regs_2_lpi_2[81:80]) , (regs_regs_2_lpi_2[83:82])
      , (regs_regs_2_lpi_2[85:84]) , (regs_regs_2_lpi_2[87:86]) , (regs_regs_2_lpi_2[89:88])
      , (regs_regs_2_lpi_2[91:90]) , (regs_regs_2_lpi_2[93:92]) , (regs_regs_2_lpi_2[95:94])
      , (regs_regs_2_lpi_2[97:96]) , (regs_regs_2_lpi_2[99:98]) , (regs_regs_2_lpi_2[101:100])
      , (regs_regs_2_lpi_2[103:102]) , (regs_regs_2_lpi_2[105:104]) , (regs_regs_2_lpi_2[107:106])
      , (regs_regs_2_lpi_2[109:108]) , (regs_regs_2_lpi_2[111:110]) , (regs_regs_2_lpi_2[113:112])
      , (regs_regs_2_lpi_2[115:114]) , (regs_regs_2_lpi_2[117:116]) , (regs_regs_2_lpi_2[119:118])
      , (regs_regs_2_lpi_2[121:120]) , (regs_regs_2_lpi_2[123:122]) , (regs_regs_2_lpi_2[125:124])
      , (regs_regs_2_lpi_2[127:126]) , (regs_regs_2_lpi_2[129:128]) , (regs_regs_2_lpi_2[131:130])
      , (regs_regs_2_lpi_2[133:132]) , (regs_regs_2_lpi_2[135:134]) , (regs_regs_2_lpi_2[137:136])
      , (regs_regs_2_lpi_2[139:138]) , (regs_regs_2_lpi_2[141:140]) , (regs_regs_2_lpi_2[143:142])
      , (regs_regs_2_lpi_2[145:144]) , (regs_regs_2_lpi_2[147:146]) , (regs_regs_2_lpi_2[149:148])
      , (regs_regs_3_lpi_2[1:0]) , (regs_regs_3_lpi_2[3:2]) , (regs_regs_3_lpi_2[5:4])
      , (regs_regs_3_lpi_2[7:6]) , (regs_regs_3_lpi_2[9:8]) , (regs_regs_3_lpi_2[11:10])
      , (regs_regs_3_lpi_2[13:12]) , (regs_regs_3_lpi_2[15:14]) , (regs_regs_3_lpi_2[17:16])
      , (regs_regs_3_lpi_2[19:18]) , (regs_regs_3_lpi_2[21:20]) , (regs_regs_3_lpi_2[23:22])
      , (regs_regs_3_lpi_2[25:24]) , (regs_regs_3_lpi_2[27:26]) , (regs_regs_3_lpi_2[29:28])
      , (regs_regs_3_lpi_2[31:30]) , (regs_regs_3_lpi_2[33:32]) , (regs_regs_3_lpi_2[35:34])
      , (regs_regs_3_lpi_2[37:36]) , (regs_regs_3_lpi_2[39:38]) , (regs_regs_3_lpi_2[41:40])
      , (regs_regs_3_lpi_2[43:42]) , (regs_regs_3_lpi_2[45:44]) , (regs_regs_3_lpi_2[47:46])
      , (regs_regs_3_lpi_2[49:48]) , (regs_regs_3_lpi_2[51:50]) , (regs_regs_3_lpi_2[53:52])
      , (regs_regs_3_lpi_2[55:54]) , (regs_regs_3_lpi_2[57:56]) , (regs_regs_3_lpi_2[59:58])
      , (regs_regs_3_lpi_2[61:60]) , (regs_regs_3_lpi_2[63:62]) , (regs_regs_3_lpi_2[65:64])
      , (regs_regs_3_lpi_2[67:66]) , (regs_regs_3_lpi_2[69:68]) , (regs_regs_3_lpi_2[71:70])
      , (regs_regs_3_lpi_2[73:72]) , (regs_regs_3_lpi_2[75:74]) , (regs_regs_3_lpi_2[77:76])
      , (regs_regs_3_lpi_2[79:78]) , (regs_regs_3_lpi_2[81:80]) , (regs_regs_3_lpi_2[83:82])
      , (regs_regs_3_lpi_2[85:84]) , (regs_regs_3_lpi_2[87:86]) , (regs_regs_3_lpi_2[89:88])
      , (regs_regs_3_lpi_2[91:90]) , (regs_regs_3_lpi_2[93:92]) , (regs_regs_3_lpi_2[95:94])
      , (regs_regs_3_lpi_2[97:96]) , (regs_regs_3_lpi_2[99:98]) , (regs_regs_3_lpi_2[101:100])
      , (regs_regs_3_lpi_2[103:102]) , (regs_regs_3_lpi_2[105:104]) , (regs_regs_3_lpi_2[107:106])
      , (regs_regs_3_lpi_2[109:108]) , (regs_regs_3_lpi_2[111:110]) , (regs_regs_3_lpi_2[113:112])
      , (regs_regs_3_lpi_2[115:114]) , (regs_regs_3_lpi_2[117:116]) , (regs_regs_3_lpi_2[119:118])
      , (regs_regs_3_lpi_2[121:120]) , (regs_regs_3_lpi_2[123:122]) , (regs_regs_3_lpi_2[125:124])
      , (regs_regs_3_lpi_2[127:126]) , (regs_regs_3_lpi_2[129:128]) , (regs_regs_3_lpi_2[131:130])
      , (regs_regs_3_lpi_2[133:132]) , (regs_regs_3_lpi_2[135:134]) , (regs_regs_3_lpi_2[137:136])
      , (regs_regs_3_lpi_2[139:138]) , (regs_regs_3_lpi_2[141:140]) , (regs_regs_3_lpi_2[143:142])
      , (regs_regs_3_lpi_2[145:144]) , (regs_regs_3_lpi_2[147:146]) , (regs_regs_3_lpi_2[149:148])
      , (regs_regs_4_lpi_2[1:0]) , (regs_regs_4_lpi_2[3:2]) , (regs_regs_4_lpi_2[5:4])
      , (regs_regs_4_lpi_2[7:6]) , (regs_regs_4_lpi_2[9:8]) , (regs_regs_4_lpi_2[11:10])
      , (regs_regs_4_lpi_2[13:12]) , (regs_regs_4_lpi_2[15:14]) , (regs_regs_4_lpi_2[17:16])
      , (regs_regs_4_lpi_2[19:18]) , (regs_regs_4_lpi_2[21:20]) , (regs_regs_4_lpi_2[23:22])
      , (regs_regs_4_lpi_2[25:24]) , (regs_regs_4_lpi_2[27:26]) , (regs_regs_4_lpi_2[29:28])
      , (regs_regs_4_lpi_2[31:30]) , (regs_regs_4_lpi_2[33:32]) , (regs_regs_4_lpi_2[35:34])
      , (regs_regs_4_lpi_2[37:36]) , (regs_regs_4_lpi_2[39:38]) , (regs_regs_4_lpi_2[41:40])
      , (regs_regs_4_lpi_2[43:42]) , (regs_regs_4_lpi_2[45:44]) , (regs_regs_4_lpi_2[47:46])
      , (regs_regs_4_lpi_2[49:48]) , (regs_regs_4_lpi_2[51:50]) , (regs_regs_4_lpi_2[53:52])
      , (regs_regs_4_lpi_2[55:54]) , (regs_regs_4_lpi_2[57:56]) , (regs_regs_4_lpi_2[59:58])
      , (regs_regs_4_lpi_2[61:60]) , (regs_regs_4_lpi_2[63:62]) , (regs_regs_4_lpi_2[65:64])
      , (regs_regs_4_lpi_2[67:66]) , (regs_regs_4_lpi_2[69:68]) , (regs_regs_4_lpi_2[71:70])
      , (regs_regs_4_lpi_2[73:72]) , (regs_regs_4_lpi_2[75:74]) , (regs_regs_4_lpi_2[77:76])
      , (regs_regs_4_lpi_2[79:78]) , (regs_regs_4_lpi_2[81:80]) , (regs_regs_4_lpi_2[83:82])
      , (regs_regs_4_lpi_2[85:84]) , (regs_regs_4_lpi_2[87:86]) , (regs_regs_4_lpi_2[89:88])
      , (regs_regs_4_lpi_2[91:90]) , (regs_regs_4_lpi_2[93:92]) , (regs_regs_4_lpi_2[95:94])
      , (regs_regs_4_lpi_2[97:96]) , (regs_regs_4_lpi_2[99:98]) , (regs_regs_4_lpi_2[101:100])
      , (regs_regs_4_lpi_2[103:102]) , (regs_regs_4_lpi_2[105:104]) , (regs_regs_4_lpi_2[107:106])
      , (regs_regs_4_lpi_2[109:108]) , (regs_regs_4_lpi_2[111:110]) , (regs_regs_4_lpi_2[113:112])
      , (regs_regs_4_lpi_2[115:114]) , (regs_regs_4_lpi_2[117:116]) , (regs_regs_4_lpi_2[119:118])
      , (regs_regs_4_lpi_2[121:120]) , (regs_regs_4_lpi_2[123:122]) , (regs_regs_4_lpi_2[125:124])
      , (regs_regs_4_lpi_2[127:126]) , (regs_regs_4_lpi_2[129:128]) , (regs_regs_4_lpi_2[131:130])
      , (regs_regs_4_lpi_2[133:132]) , (regs_regs_4_lpi_2[135:134]) , (regs_regs_4_lpi_2[137:136])
      , (regs_regs_4_lpi_2[139:138]) , (regs_regs_4_lpi_2[141:140]) , (regs_regs_4_lpi_2[143:142])
      , (regs_regs_4_lpi_2[145:144]) , (regs_regs_4_lpi_2[147:146]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg12 = MUX_v_2_512_2({(regs_regs_0_lpi_2[25:24]) , (regs_regs_0_lpi_2[27:26])
      , (regs_regs_0_lpi_2[29:28]) , (regs_regs_0_lpi_2[31:30]) , (regs_regs_0_lpi_2[33:32])
      , (regs_regs_0_lpi_2[35:34]) , (regs_regs_0_lpi_2[37:36]) , (regs_regs_0_lpi_2[39:38])
      , (regs_regs_0_lpi_2[41:40]) , (regs_regs_0_lpi_2[43:42]) , (regs_regs_0_lpi_2[45:44])
      , (regs_regs_0_lpi_2[47:46]) , (regs_regs_0_lpi_2[49:48]) , (regs_regs_0_lpi_2[51:50])
      , (regs_regs_0_lpi_2[53:52]) , (regs_regs_0_lpi_2[55:54]) , (regs_regs_0_lpi_2[57:56])
      , (regs_regs_0_lpi_2[59:58]) , (regs_regs_0_lpi_2[61:60]) , (regs_regs_0_lpi_2[63:62])
      , (regs_regs_0_lpi_2[65:64]) , (regs_regs_0_lpi_2[67:66]) , (regs_regs_0_lpi_2[69:68])
      , (regs_regs_0_lpi_2[71:70]) , (regs_regs_0_lpi_2[73:72]) , (regs_regs_0_lpi_2[75:74])
      , (regs_regs_0_lpi_2[77:76]) , (regs_regs_0_lpi_2[79:78]) , (regs_regs_0_lpi_2[81:80])
      , (regs_regs_0_lpi_2[83:82]) , (regs_regs_0_lpi_2[85:84]) , (regs_regs_0_lpi_2[87:86])
      , (regs_regs_0_lpi_2[89:88]) , (regs_regs_0_lpi_2[91:90]) , (regs_regs_0_lpi_2[93:92])
      , (regs_regs_0_lpi_2[95:94]) , (regs_regs_0_lpi_2[97:96]) , (regs_regs_0_lpi_2[99:98])
      , (regs_regs_0_lpi_2[101:100]) , (regs_regs_0_lpi_2[103:102]) , (regs_regs_0_lpi_2[105:104])
      , (regs_regs_0_lpi_2[107:106]) , (regs_regs_0_lpi_2[109:108]) , (regs_regs_0_lpi_2[111:110])
      , (regs_regs_0_lpi_2[113:112]) , (regs_regs_0_lpi_2[115:114]) , (regs_regs_0_lpi_2[117:116])
      , (regs_regs_0_lpi_2[119:118]) , (regs_regs_0_lpi_2[121:120]) , (regs_regs_0_lpi_2[123:122])
      , (regs_regs_0_lpi_2[125:124]) , (regs_regs_0_lpi_2[127:126]) , (regs_regs_0_lpi_2[129:128])
      , (regs_regs_0_lpi_2[131:130]) , (regs_regs_0_lpi_2[133:132]) , (regs_regs_0_lpi_2[135:134])
      , (regs_regs_0_lpi_2[137:136]) , (regs_regs_0_lpi_2[139:138]) , (regs_regs_0_lpi_2[141:140])
      , (regs_regs_0_lpi_2[143:142]) , (regs_regs_0_lpi_2[145:144]) , (regs_regs_0_lpi_2[147:146])
      , (regs_regs_0_lpi_2[149:148]) , (regs_regs_1_lpi_2[1:0]) , (regs_regs_1_lpi_2[3:2])
      , (regs_regs_1_lpi_2[5:4]) , (regs_regs_1_lpi_2[7:6]) , (regs_regs_1_lpi_2[9:8])
      , (regs_regs_1_lpi_2[11:10]) , (regs_regs_1_lpi_2[13:12]) , (regs_regs_1_lpi_2[15:14])
      , (regs_regs_1_lpi_2[17:16]) , (regs_regs_1_lpi_2[19:18]) , (regs_regs_1_lpi_2[21:20])
      , (regs_regs_1_lpi_2[23:22]) , (regs_regs_1_lpi_2[25:24]) , (regs_regs_1_lpi_2[27:26])
      , (regs_regs_1_lpi_2[29:28]) , (regs_regs_1_lpi_2[31:30]) , (regs_regs_1_lpi_2[33:32])
      , (regs_regs_1_lpi_2[35:34]) , (regs_regs_1_lpi_2[37:36]) , (regs_regs_1_lpi_2[39:38])
      , (regs_regs_1_lpi_2[41:40]) , (regs_regs_1_lpi_2[43:42]) , (regs_regs_1_lpi_2[45:44])
      , (regs_regs_1_lpi_2[47:46]) , (regs_regs_1_lpi_2[49:48]) , (regs_regs_1_lpi_2[51:50])
      , (regs_regs_1_lpi_2[53:52]) , (regs_regs_1_lpi_2[55:54]) , (regs_regs_1_lpi_2[57:56])
      , (regs_regs_1_lpi_2[59:58]) , (regs_regs_1_lpi_2[61:60]) , (regs_regs_1_lpi_2[63:62])
      , (regs_regs_1_lpi_2[65:64]) , (regs_regs_1_lpi_2[67:66]) , (regs_regs_1_lpi_2[69:68])
      , (regs_regs_1_lpi_2[71:70]) , (regs_regs_1_lpi_2[73:72]) , (regs_regs_1_lpi_2[75:74])
      , (regs_regs_1_lpi_2[77:76]) , (regs_regs_1_lpi_2[79:78]) , (regs_regs_1_lpi_2[81:80])
      , (regs_regs_1_lpi_2[83:82]) , (regs_regs_1_lpi_2[85:84]) , (regs_regs_1_lpi_2[87:86])
      , (regs_regs_1_lpi_2[89:88]) , (regs_regs_1_lpi_2[91:90]) , (regs_regs_1_lpi_2[93:92])
      , (regs_regs_1_lpi_2[95:94]) , (regs_regs_1_lpi_2[97:96]) , (regs_regs_1_lpi_2[99:98])
      , (regs_regs_1_lpi_2[101:100]) , (regs_regs_1_lpi_2[103:102]) , (regs_regs_1_lpi_2[105:104])
      , (regs_regs_1_lpi_2[107:106]) , (regs_regs_1_lpi_2[109:108]) , (regs_regs_1_lpi_2[111:110])
      , (regs_regs_1_lpi_2[113:112]) , (regs_regs_1_lpi_2[115:114]) , (regs_regs_1_lpi_2[117:116])
      , (regs_regs_1_lpi_2[119:118]) , (regs_regs_1_lpi_2[121:120]) , (regs_regs_1_lpi_2[123:122])
      , (regs_regs_1_lpi_2[125:124]) , (regs_regs_1_lpi_2[127:126]) , (regs_regs_1_lpi_2[129:128])
      , (regs_regs_1_lpi_2[131:130]) , (regs_regs_1_lpi_2[133:132]) , (regs_regs_1_lpi_2[135:134])
      , (regs_regs_1_lpi_2[137:136]) , (regs_regs_1_lpi_2[139:138]) , (regs_regs_1_lpi_2[141:140])
      , (regs_regs_1_lpi_2[143:142]) , (regs_regs_1_lpi_2[145:144]) , (regs_regs_1_lpi_2[147:146])
      , (regs_regs_1_lpi_2[149:148]) , (regs_regs_2_lpi_2[1:0]) , (regs_regs_2_lpi_2[3:2])
      , (regs_regs_2_lpi_2[5:4]) , (regs_regs_2_lpi_2[7:6]) , (regs_regs_2_lpi_2[9:8])
      , (regs_regs_2_lpi_2[11:10]) , (regs_regs_2_lpi_2[13:12]) , (regs_regs_2_lpi_2[15:14])
      , (regs_regs_2_lpi_2[17:16]) , (regs_regs_2_lpi_2[19:18]) , (regs_regs_2_lpi_2[21:20])
      , (regs_regs_2_lpi_2[23:22]) , (regs_regs_2_lpi_2[25:24]) , (regs_regs_2_lpi_2[27:26])
      , (regs_regs_2_lpi_2[29:28]) , (regs_regs_2_lpi_2[31:30]) , (regs_regs_2_lpi_2[33:32])
      , (regs_regs_2_lpi_2[35:34]) , (regs_regs_2_lpi_2[37:36]) , (regs_regs_2_lpi_2[39:38])
      , (regs_regs_2_lpi_2[41:40]) , (regs_regs_2_lpi_2[43:42]) , (regs_regs_2_lpi_2[45:44])
      , (regs_regs_2_lpi_2[47:46]) , (regs_regs_2_lpi_2[49:48]) , (regs_regs_2_lpi_2[51:50])
      , (regs_regs_2_lpi_2[53:52]) , (regs_regs_2_lpi_2[55:54]) , (regs_regs_2_lpi_2[57:56])
      , (regs_regs_2_lpi_2[59:58]) , (regs_regs_2_lpi_2[61:60]) , (regs_regs_2_lpi_2[63:62])
      , (regs_regs_2_lpi_2[65:64]) , (regs_regs_2_lpi_2[67:66]) , (regs_regs_2_lpi_2[69:68])
      , (regs_regs_2_lpi_2[71:70]) , (regs_regs_2_lpi_2[73:72]) , (regs_regs_2_lpi_2[75:74])
      , (regs_regs_2_lpi_2[77:76]) , (regs_regs_2_lpi_2[79:78]) , (regs_regs_2_lpi_2[81:80])
      , (regs_regs_2_lpi_2[83:82]) , (regs_regs_2_lpi_2[85:84]) , (regs_regs_2_lpi_2[87:86])
      , (regs_regs_2_lpi_2[89:88]) , (regs_regs_2_lpi_2[91:90]) , (regs_regs_2_lpi_2[93:92])
      , (regs_regs_2_lpi_2[95:94]) , (regs_regs_2_lpi_2[97:96]) , (regs_regs_2_lpi_2[99:98])
      , (regs_regs_2_lpi_2[101:100]) , (regs_regs_2_lpi_2[103:102]) , (regs_regs_2_lpi_2[105:104])
      , (regs_regs_2_lpi_2[107:106]) , (regs_regs_2_lpi_2[109:108]) , (regs_regs_2_lpi_2[111:110])
      , (regs_regs_2_lpi_2[113:112]) , (regs_regs_2_lpi_2[115:114]) , (regs_regs_2_lpi_2[117:116])
      , (regs_regs_2_lpi_2[119:118]) , (regs_regs_2_lpi_2[121:120]) , (regs_regs_2_lpi_2[123:122])
      , (regs_regs_2_lpi_2[125:124]) , (regs_regs_2_lpi_2[127:126]) , (regs_regs_2_lpi_2[129:128])
      , (regs_regs_2_lpi_2[131:130]) , (regs_regs_2_lpi_2[133:132]) , (regs_regs_2_lpi_2[135:134])
      , (regs_regs_2_lpi_2[137:136]) , (regs_regs_2_lpi_2[139:138]) , (regs_regs_2_lpi_2[141:140])
      , (regs_regs_2_lpi_2[143:142]) , (regs_regs_2_lpi_2[145:144]) , (regs_regs_2_lpi_2[147:146])
      , (regs_regs_2_lpi_2[149:148]) , (regs_regs_3_lpi_2[1:0]) , (regs_regs_3_lpi_2[3:2])
      , (regs_regs_3_lpi_2[5:4]) , (regs_regs_3_lpi_2[7:6]) , (regs_regs_3_lpi_2[9:8])
      , (regs_regs_3_lpi_2[11:10]) , (regs_regs_3_lpi_2[13:12]) , (regs_regs_3_lpi_2[15:14])
      , (regs_regs_3_lpi_2[17:16]) , (regs_regs_3_lpi_2[19:18]) , (regs_regs_3_lpi_2[21:20])
      , (regs_regs_3_lpi_2[23:22]) , (regs_regs_3_lpi_2[25:24]) , (regs_regs_3_lpi_2[27:26])
      , (regs_regs_3_lpi_2[29:28]) , (regs_regs_3_lpi_2[31:30]) , (regs_regs_3_lpi_2[33:32])
      , (regs_regs_3_lpi_2[35:34]) , (regs_regs_3_lpi_2[37:36]) , (regs_regs_3_lpi_2[39:38])
      , (regs_regs_3_lpi_2[41:40]) , (regs_regs_3_lpi_2[43:42]) , (regs_regs_3_lpi_2[45:44])
      , (regs_regs_3_lpi_2[47:46]) , (regs_regs_3_lpi_2[49:48]) , (regs_regs_3_lpi_2[51:50])
      , (regs_regs_3_lpi_2[53:52]) , (regs_regs_3_lpi_2[55:54]) , (regs_regs_3_lpi_2[57:56])
      , (regs_regs_3_lpi_2[59:58]) , (regs_regs_3_lpi_2[61:60]) , (regs_regs_3_lpi_2[63:62])
      , (regs_regs_3_lpi_2[65:64]) , (regs_regs_3_lpi_2[67:66]) , (regs_regs_3_lpi_2[69:68])
      , (regs_regs_3_lpi_2[71:70]) , (regs_regs_3_lpi_2[73:72]) , (regs_regs_3_lpi_2[75:74])
      , (regs_regs_3_lpi_2[77:76]) , (regs_regs_3_lpi_2[79:78]) , (regs_regs_3_lpi_2[81:80])
      , (regs_regs_3_lpi_2[83:82]) , (regs_regs_3_lpi_2[85:84]) , (regs_regs_3_lpi_2[87:86])
      , (regs_regs_3_lpi_2[89:88]) , (regs_regs_3_lpi_2[91:90]) , (regs_regs_3_lpi_2[93:92])
      , (regs_regs_3_lpi_2[95:94]) , (regs_regs_3_lpi_2[97:96]) , (regs_regs_3_lpi_2[99:98])
      , (regs_regs_3_lpi_2[101:100]) , (regs_regs_3_lpi_2[103:102]) , (regs_regs_3_lpi_2[105:104])
      , (regs_regs_3_lpi_2[107:106]) , (regs_regs_3_lpi_2[109:108]) , (regs_regs_3_lpi_2[111:110])
      , (regs_regs_3_lpi_2[113:112]) , (regs_regs_3_lpi_2[115:114]) , (regs_regs_3_lpi_2[117:116])
      , (regs_regs_3_lpi_2[119:118]) , (regs_regs_3_lpi_2[121:120]) , (regs_regs_3_lpi_2[123:122])
      , (regs_regs_3_lpi_2[125:124]) , (regs_regs_3_lpi_2[127:126]) , (regs_regs_3_lpi_2[129:128])
      , (regs_regs_3_lpi_2[131:130]) , (regs_regs_3_lpi_2[133:132]) , (regs_regs_3_lpi_2[135:134])
      , (regs_regs_3_lpi_2[137:136]) , (regs_regs_3_lpi_2[139:138]) , (regs_regs_3_lpi_2[141:140])
      , (regs_regs_3_lpi_2[143:142]) , (regs_regs_3_lpi_2[145:144]) , (regs_regs_3_lpi_2[147:146])
      , (regs_regs_3_lpi_2[149:148]) , (regs_regs_4_lpi_2[1:0]) , (regs_regs_4_lpi_2[3:2])
      , (regs_regs_4_lpi_2[5:4]) , (regs_regs_4_lpi_2[7:6]) , (regs_regs_4_lpi_2[9:8])
      , (regs_regs_4_lpi_2[11:10]) , (regs_regs_4_lpi_2[13:12]) , (regs_regs_4_lpi_2[15:14])
      , (regs_regs_4_lpi_2[17:16]) , (regs_regs_4_lpi_2[19:18]) , (regs_regs_4_lpi_2[21:20])
      , (regs_regs_4_lpi_2[23:22]) , (regs_regs_4_lpi_2[25:24]) , (regs_regs_4_lpi_2[27:26])
      , (regs_regs_4_lpi_2[29:28]) , (regs_regs_4_lpi_2[31:30]) , (regs_regs_4_lpi_2[33:32])
      , (regs_regs_4_lpi_2[35:34]) , (regs_regs_4_lpi_2[37:36]) , (regs_regs_4_lpi_2[39:38])
      , (regs_regs_4_lpi_2[41:40]) , (regs_regs_4_lpi_2[43:42]) , (regs_regs_4_lpi_2[45:44])
      , (regs_regs_4_lpi_2[47:46]) , (regs_regs_4_lpi_2[49:48]) , (regs_regs_4_lpi_2[51:50])
      , (regs_regs_4_lpi_2[53:52]) , (regs_regs_4_lpi_2[55:54]) , (regs_regs_4_lpi_2[57:56])
      , (regs_regs_4_lpi_2[59:58]) , (regs_regs_4_lpi_2[61:60]) , (regs_regs_4_lpi_2[63:62])
      , (regs_regs_4_lpi_2[65:64]) , (regs_regs_4_lpi_2[67:66]) , (regs_regs_4_lpi_2[69:68])
      , (regs_regs_4_lpi_2[71:70]) , (regs_regs_4_lpi_2[73:72]) , (regs_regs_4_lpi_2[75:74])
      , (regs_regs_4_lpi_2[77:76]) , (regs_regs_4_lpi_2[79:78]) , (regs_regs_4_lpi_2[81:80])
      , (regs_regs_4_lpi_2[83:82]) , (regs_regs_4_lpi_2[85:84]) , (regs_regs_4_lpi_2[87:86])
      , (regs_regs_4_lpi_2[89:88]) , (regs_regs_4_lpi_2[91:90]) , (regs_regs_4_lpi_2[93:92])
      , (regs_regs_4_lpi_2[95:94]) , (regs_regs_4_lpi_2[97:96]) , (regs_regs_4_lpi_2[99:98])
      , (regs_regs_4_lpi_2[101:100]) , (regs_regs_4_lpi_2[103:102]) , (regs_regs_4_lpi_2[105:104])
      , (regs_regs_4_lpi_2[107:106]) , (regs_regs_4_lpi_2[109:108]) , (regs_regs_4_lpi_2[111:110])
      , (regs_regs_4_lpi_2[113:112]) , (regs_regs_4_lpi_2[115:114]) , (regs_regs_4_lpi_2[117:116])
      , (regs_regs_4_lpi_2[119:118]) , (regs_regs_4_lpi_2[121:120]) , (regs_regs_4_lpi_2[123:122])
      , (regs_regs_4_lpi_2[125:124]) , (regs_regs_4_lpi_2[127:126]) , (regs_regs_4_lpi_2[129:128])
      , (regs_regs_4_lpi_2[131:130]) , (regs_regs_4_lpi_2[133:132]) , (regs_regs_4_lpi_2[135:134])
      , (regs_regs_4_lpi_2[137:136]) , (regs_regs_4_lpi_2[139:138]) , (regs_regs_4_lpi_2[141:140])
      , (regs_regs_4_lpi_2[143:142]) , (regs_regs_4_lpi_2[145:144]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg11 = MUX_v_2_512_2({(regs_regs_0_lpi_2[23:22]) , (regs_regs_0_lpi_2[25:24])
      , (regs_regs_0_lpi_2[27:26]) , (regs_regs_0_lpi_2[29:28]) , (regs_regs_0_lpi_2[31:30])
      , (regs_regs_0_lpi_2[33:32]) , (regs_regs_0_lpi_2[35:34]) , (regs_regs_0_lpi_2[37:36])
      , (regs_regs_0_lpi_2[39:38]) , (regs_regs_0_lpi_2[41:40]) , (regs_regs_0_lpi_2[43:42])
      , (regs_regs_0_lpi_2[45:44]) , (regs_regs_0_lpi_2[47:46]) , (regs_regs_0_lpi_2[49:48])
      , (regs_regs_0_lpi_2[51:50]) , (regs_regs_0_lpi_2[53:52]) , (regs_regs_0_lpi_2[55:54])
      , (regs_regs_0_lpi_2[57:56]) , (regs_regs_0_lpi_2[59:58]) , (regs_regs_0_lpi_2[61:60])
      , (regs_regs_0_lpi_2[63:62]) , (regs_regs_0_lpi_2[65:64]) , (regs_regs_0_lpi_2[67:66])
      , (regs_regs_0_lpi_2[69:68]) , (regs_regs_0_lpi_2[71:70]) , (regs_regs_0_lpi_2[73:72])
      , (regs_regs_0_lpi_2[75:74]) , (regs_regs_0_lpi_2[77:76]) , (regs_regs_0_lpi_2[79:78])
      , (regs_regs_0_lpi_2[81:80]) , (regs_regs_0_lpi_2[83:82]) , (regs_regs_0_lpi_2[85:84])
      , (regs_regs_0_lpi_2[87:86]) , (regs_regs_0_lpi_2[89:88]) , (regs_regs_0_lpi_2[91:90])
      , (regs_regs_0_lpi_2[93:92]) , (regs_regs_0_lpi_2[95:94]) , (regs_regs_0_lpi_2[97:96])
      , (regs_regs_0_lpi_2[99:98]) , (regs_regs_0_lpi_2[101:100]) , (regs_regs_0_lpi_2[103:102])
      , (regs_regs_0_lpi_2[105:104]) , (regs_regs_0_lpi_2[107:106]) , (regs_regs_0_lpi_2[109:108])
      , (regs_regs_0_lpi_2[111:110]) , (regs_regs_0_lpi_2[113:112]) , (regs_regs_0_lpi_2[115:114])
      , (regs_regs_0_lpi_2[117:116]) , (regs_regs_0_lpi_2[119:118]) , (regs_regs_0_lpi_2[121:120])
      , (regs_regs_0_lpi_2[123:122]) , (regs_regs_0_lpi_2[125:124]) , (regs_regs_0_lpi_2[127:126])
      , (regs_regs_0_lpi_2[129:128]) , (regs_regs_0_lpi_2[131:130]) , (regs_regs_0_lpi_2[133:132])
      , (regs_regs_0_lpi_2[135:134]) , (regs_regs_0_lpi_2[137:136]) , (regs_regs_0_lpi_2[139:138])
      , (regs_regs_0_lpi_2[141:140]) , (regs_regs_0_lpi_2[143:142]) , (regs_regs_0_lpi_2[145:144])
      , (regs_regs_0_lpi_2[147:146]) , (regs_regs_0_lpi_2[149:148]) , (regs_regs_1_lpi_2[1:0])
      , (regs_regs_1_lpi_2[3:2]) , (regs_regs_1_lpi_2[5:4]) , (regs_regs_1_lpi_2[7:6])
      , (regs_regs_1_lpi_2[9:8]) , (regs_regs_1_lpi_2[11:10]) , (regs_regs_1_lpi_2[13:12])
      , (regs_regs_1_lpi_2[15:14]) , (regs_regs_1_lpi_2[17:16]) , (regs_regs_1_lpi_2[19:18])
      , (regs_regs_1_lpi_2[21:20]) , (regs_regs_1_lpi_2[23:22]) , (regs_regs_1_lpi_2[25:24])
      , (regs_regs_1_lpi_2[27:26]) , (regs_regs_1_lpi_2[29:28]) , (regs_regs_1_lpi_2[31:30])
      , (regs_regs_1_lpi_2[33:32]) , (regs_regs_1_lpi_2[35:34]) , (regs_regs_1_lpi_2[37:36])
      , (regs_regs_1_lpi_2[39:38]) , (regs_regs_1_lpi_2[41:40]) , (regs_regs_1_lpi_2[43:42])
      , (regs_regs_1_lpi_2[45:44]) , (regs_regs_1_lpi_2[47:46]) , (regs_regs_1_lpi_2[49:48])
      , (regs_regs_1_lpi_2[51:50]) , (regs_regs_1_lpi_2[53:52]) , (regs_regs_1_lpi_2[55:54])
      , (regs_regs_1_lpi_2[57:56]) , (regs_regs_1_lpi_2[59:58]) , (regs_regs_1_lpi_2[61:60])
      , (regs_regs_1_lpi_2[63:62]) , (regs_regs_1_lpi_2[65:64]) , (regs_regs_1_lpi_2[67:66])
      , (regs_regs_1_lpi_2[69:68]) , (regs_regs_1_lpi_2[71:70]) , (regs_regs_1_lpi_2[73:72])
      , (regs_regs_1_lpi_2[75:74]) , (regs_regs_1_lpi_2[77:76]) , (regs_regs_1_lpi_2[79:78])
      , (regs_regs_1_lpi_2[81:80]) , (regs_regs_1_lpi_2[83:82]) , (regs_regs_1_lpi_2[85:84])
      , (regs_regs_1_lpi_2[87:86]) , (regs_regs_1_lpi_2[89:88]) , (regs_regs_1_lpi_2[91:90])
      , (regs_regs_1_lpi_2[93:92]) , (regs_regs_1_lpi_2[95:94]) , (regs_regs_1_lpi_2[97:96])
      , (regs_regs_1_lpi_2[99:98]) , (regs_regs_1_lpi_2[101:100]) , (regs_regs_1_lpi_2[103:102])
      , (regs_regs_1_lpi_2[105:104]) , (regs_regs_1_lpi_2[107:106]) , (regs_regs_1_lpi_2[109:108])
      , (regs_regs_1_lpi_2[111:110]) , (regs_regs_1_lpi_2[113:112]) , (regs_regs_1_lpi_2[115:114])
      , (regs_regs_1_lpi_2[117:116]) , (regs_regs_1_lpi_2[119:118]) , (regs_regs_1_lpi_2[121:120])
      , (regs_regs_1_lpi_2[123:122]) , (regs_regs_1_lpi_2[125:124]) , (regs_regs_1_lpi_2[127:126])
      , (regs_regs_1_lpi_2[129:128]) , (regs_regs_1_lpi_2[131:130]) , (regs_regs_1_lpi_2[133:132])
      , (regs_regs_1_lpi_2[135:134]) , (regs_regs_1_lpi_2[137:136]) , (regs_regs_1_lpi_2[139:138])
      , (regs_regs_1_lpi_2[141:140]) , (regs_regs_1_lpi_2[143:142]) , (regs_regs_1_lpi_2[145:144])
      , (regs_regs_1_lpi_2[147:146]) , (regs_regs_1_lpi_2[149:148]) , (regs_regs_2_lpi_2[1:0])
      , (regs_regs_2_lpi_2[3:2]) , (regs_regs_2_lpi_2[5:4]) , (regs_regs_2_lpi_2[7:6])
      , (regs_regs_2_lpi_2[9:8]) , (regs_regs_2_lpi_2[11:10]) , (regs_regs_2_lpi_2[13:12])
      , (regs_regs_2_lpi_2[15:14]) , (regs_regs_2_lpi_2[17:16]) , (regs_regs_2_lpi_2[19:18])
      , (regs_regs_2_lpi_2[21:20]) , (regs_regs_2_lpi_2[23:22]) , (regs_regs_2_lpi_2[25:24])
      , (regs_regs_2_lpi_2[27:26]) , (regs_regs_2_lpi_2[29:28]) , (regs_regs_2_lpi_2[31:30])
      , (regs_regs_2_lpi_2[33:32]) , (regs_regs_2_lpi_2[35:34]) , (regs_regs_2_lpi_2[37:36])
      , (regs_regs_2_lpi_2[39:38]) , (regs_regs_2_lpi_2[41:40]) , (regs_regs_2_lpi_2[43:42])
      , (regs_regs_2_lpi_2[45:44]) , (regs_regs_2_lpi_2[47:46]) , (regs_regs_2_lpi_2[49:48])
      , (regs_regs_2_lpi_2[51:50]) , (regs_regs_2_lpi_2[53:52]) , (regs_regs_2_lpi_2[55:54])
      , (regs_regs_2_lpi_2[57:56]) , (regs_regs_2_lpi_2[59:58]) , (regs_regs_2_lpi_2[61:60])
      , (regs_regs_2_lpi_2[63:62]) , (regs_regs_2_lpi_2[65:64]) , (regs_regs_2_lpi_2[67:66])
      , (regs_regs_2_lpi_2[69:68]) , (regs_regs_2_lpi_2[71:70]) , (regs_regs_2_lpi_2[73:72])
      , (regs_regs_2_lpi_2[75:74]) , (regs_regs_2_lpi_2[77:76]) , (regs_regs_2_lpi_2[79:78])
      , (regs_regs_2_lpi_2[81:80]) , (regs_regs_2_lpi_2[83:82]) , (regs_regs_2_lpi_2[85:84])
      , (regs_regs_2_lpi_2[87:86]) , (regs_regs_2_lpi_2[89:88]) , (regs_regs_2_lpi_2[91:90])
      , (regs_regs_2_lpi_2[93:92]) , (regs_regs_2_lpi_2[95:94]) , (regs_regs_2_lpi_2[97:96])
      , (regs_regs_2_lpi_2[99:98]) , (regs_regs_2_lpi_2[101:100]) , (regs_regs_2_lpi_2[103:102])
      , (regs_regs_2_lpi_2[105:104]) , (regs_regs_2_lpi_2[107:106]) , (regs_regs_2_lpi_2[109:108])
      , (regs_regs_2_lpi_2[111:110]) , (regs_regs_2_lpi_2[113:112]) , (regs_regs_2_lpi_2[115:114])
      , (regs_regs_2_lpi_2[117:116]) , (regs_regs_2_lpi_2[119:118]) , (regs_regs_2_lpi_2[121:120])
      , (regs_regs_2_lpi_2[123:122]) , (regs_regs_2_lpi_2[125:124]) , (regs_regs_2_lpi_2[127:126])
      , (regs_regs_2_lpi_2[129:128]) , (regs_regs_2_lpi_2[131:130]) , (regs_regs_2_lpi_2[133:132])
      , (regs_regs_2_lpi_2[135:134]) , (regs_regs_2_lpi_2[137:136]) , (regs_regs_2_lpi_2[139:138])
      , (regs_regs_2_lpi_2[141:140]) , (regs_regs_2_lpi_2[143:142]) , (regs_regs_2_lpi_2[145:144])
      , (regs_regs_2_lpi_2[147:146]) , (regs_regs_2_lpi_2[149:148]) , (regs_regs_3_lpi_2[1:0])
      , (regs_regs_3_lpi_2[3:2]) , (regs_regs_3_lpi_2[5:4]) , (regs_regs_3_lpi_2[7:6])
      , (regs_regs_3_lpi_2[9:8]) , (regs_regs_3_lpi_2[11:10]) , (regs_regs_3_lpi_2[13:12])
      , (regs_regs_3_lpi_2[15:14]) , (regs_regs_3_lpi_2[17:16]) , (regs_regs_3_lpi_2[19:18])
      , (regs_regs_3_lpi_2[21:20]) , (regs_regs_3_lpi_2[23:22]) , (regs_regs_3_lpi_2[25:24])
      , (regs_regs_3_lpi_2[27:26]) , (regs_regs_3_lpi_2[29:28]) , (regs_regs_3_lpi_2[31:30])
      , (regs_regs_3_lpi_2[33:32]) , (regs_regs_3_lpi_2[35:34]) , (regs_regs_3_lpi_2[37:36])
      , (regs_regs_3_lpi_2[39:38]) , (regs_regs_3_lpi_2[41:40]) , (regs_regs_3_lpi_2[43:42])
      , (regs_regs_3_lpi_2[45:44]) , (regs_regs_3_lpi_2[47:46]) , (regs_regs_3_lpi_2[49:48])
      , (regs_regs_3_lpi_2[51:50]) , (regs_regs_3_lpi_2[53:52]) , (regs_regs_3_lpi_2[55:54])
      , (regs_regs_3_lpi_2[57:56]) , (regs_regs_3_lpi_2[59:58]) , (regs_regs_3_lpi_2[61:60])
      , (regs_regs_3_lpi_2[63:62]) , (regs_regs_3_lpi_2[65:64]) , (regs_regs_3_lpi_2[67:66])
      , (regs_regs_3_lpi_2[69:68]) , (regs_regs_3_lpi_2[71:70]) , (regs_regs_3_lpi_2[73:72])
      , (regs_regs_3_lpi_2[75:74]) , (regs_regs_3_lpi_2[77:76]) , (regs_regs_3_lpi_2[79:78])
      , (regs_regs_3_lpi_2[81:80]) , (regs_regs_3_lpi_2[83:82]) , (regs_regs_3_lpi_2[85:84])
      , (regs_regs_3_lpi_2[87:86]) , (regs_regs_3_lpi_2[89:88]) , (regs_regs_3_lpi_2[91:90])
      , (regs_regs_3_lpi_2[93:92]) , (regs_regs_3_lpi_2[95:94]) , (regs_regs_3_lpi_2[97:96])
      , (regs_regs_3_lpi_2[99:98]) , (regs_regs_3_lpi_2[101:100]) , (regs_regs_3_lpi_2[103:102])
      , (regs_regs_3_lpi_2[105:104]) , (regs_regs_3_lpi_2[107:106]) , (regs_regs_3_lpi_2[109:108])
      , (regs_regs_3_lpi_2[111:110]) , (regs_regs_3_lpi_2[113:112]) , (regs_regs_3_lpi_2[115:114])
      , (regs_regs_3_lpi_2[117:116]) , (regs_regs_3_lpi_2[119:118]) , (regs_regs_3_lpi_2[121:120])
      , (regs_regs_3_lpi_2[123:122]) , (regs_regs_3_lpi_2[125:124]) , (regs_regs_3_lpi_2[127:126])
      , (regs_regs_3_lpi_2[129:128]) , (regs_regs_3_lpi_2[131:130]) , (regs_regs_3_lpi_2[133:132])
      , (regs_regs_3_lpi_2[135:134]) , (regs_regs_3_lpi_2[137:136]) , (regs_regs_3_lpi_2[139:138])
      , (regs_regs_3_lpi_2[141:140]) , (regs_regs_3_lpi_2[143:142]) , (regs_regs_3_lpi_2[145:144])
      , (regs_regs_3_lpi_2[147:146]) , (regs_regs_3_lpi_2[149:148]) , (regs_regs_4_lpi_2[1:0])
      , (regs_regs_4_lpi_2[3:2]) , (regs_regs_4_lpi_2[5:4]) , (regs_regs_4_lpi_2[7:6])
      , (regs_regs_4_lpi_2[9:8]) , (regs_regs_4_lpi_2[11:10]) , (regs_regs_4_lpi_2[13:12])
      , (regs_regs_4_lpi_2[15:14]) , (regs_regs_4_lpi_2[17:16]) , (regs_regs_4_lpi_2[19:18])
      , (regs_regs_4_lpi_2[21:20]) , (regs_regs_4_lpi_2[23:22]) , (regs_regs_4_lpi_2[25:24])
      , (regs_regs_4_lpi_2[27:26]) , (regs_regs_4_lpi_2[29:28]) , (regs_regs_4_lpi_2[31:30])
      , (regs_regs_4_lpi_2[33:32]) , (regs_regs_4_lpi_2[35:34]) , (regs_regs_4_lpi_2[37:36])
      , (regs_regs_4_lpi_2[39:38]) , (regs_regs_4_lpi_2[41:40]) , (regs_regs_4_lpi_2[43:42])
      , (regs_regs_4_lpi_2[45:44]) , (regs_regs_4_lpi_2[47:46]) , (regs_regs_4_lpi_2[49:48])
      , (regs_regs_4_lpi_2[51:50]) , (regs_regs_4_lpi_2[53:52]) , (regs_regs_4_lpi_2[55:54])
      , (regs_regs_4_lpi_2[57:56]) , (regs_regs_4_lpi_2[59:58]) , (regs_regs_4_lpi_2[61:60])
      , (regs_regs_4_lpi_2[63:62]) , (regs_regs_4_lpi_2[65:64]) , (regs_regs_4_lpi_2[67:66])
      , (regs_regs_4_lpi_2[69:68]) , (regs_regs_4_lpi_2[71:70]) , (regs_regs_4_lpi_2[73:72])
      , (regs_regs_4_lpi_2[75:74]) , (regs_regs_4_lpi_2[77:76]) , (regs_regs_4_lpi_2[79:78])
      , (regs_regs_4_lpi_2[81:80]) , (regs_regs_4_lpi_2[83:82]) , (regs_regs_4_lpi_2[85:84])
      , (regs_regs_4_lpi_2[87:86]) , (regs_regs_4_lpi_2[89:88]) , (regs_regs_4_lpi_2[91:90])
      , (regs_regs_4_lpi_2[93:92]) , (regs_regs_4_lpi_2[95:94]) , (regs_regs_4_lpi_2[97:96])
      , (regs_regs_4_lpi_2[99:98]) , (regs_regs_4_lpi_2[101:100]) , (regs_regs_4_lpi_2[103:102])
      , (regs_regs_4_lpi_2[105:104]) , (regs_regs_4_lpi_2[107:106]) , (regs_regs_4_lpi_2[109:108])
      , (regs_regs_4_lpi_2[111:110]) , (regs_regs_4_lpi_2[113:112]) , (regs_regs_4_lpi_2[115:114])
      , (regs_regs_4_lpi_2[117:116]) , (regs_regs_4_lpi_2[119:118]) , (regs_regs_4_lpi_2[121:120])
      , (regs_regs_4_lpi_2[123:122]) , (regs_regs_4_lpi_2[125:124]) , (regs_regs_4_lpi_2[127:126])
      , (regs_regs_4_lpi_2[129:128]) , (regs_regs_4_lpi_2[131:130]) , (regs_regs_4_lpi_2[133:132])
      , (regs_regs_4_lpi_2[135:134]) , (regs_regs_4_lpi_2[137:136]) , (regs_regs_4_lpi_2[139:138])
      , (regs_regs_4_lpi_2[141:140]) , (regs_regs_4_lpi_2[143:142]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg10 = MUX_v_2_512_2({(regs_regs_0_lpi_2[21:20]) , (regs_regs_0_lpi_2[23:22])
      , (regs_regs_0_lpi_2[25:24]) , (regs_regs_0_lpi_2[27:26]) , (regs_regs_0_lpi_2[29:28])
      , (regs_regs_0_lpi_2[31:30]) , (regs_regs_0_lpi_2[33:32]) , (regs_regs_0_lpi_2[35:34])
      , (regs_regs_0_lpi_2[37:36]) , (regs_regs_0_lpi_2[39:38]) , (regs_regs_0_lpi_2[41:40])
      , (regs_regs_0_lpi_2[43:42]) , (regs_regs_0_lpi_2[45:44]) , (regs_regs_0_lpi_2[47:46])
      , (regs_regs_0_lpi_2[49:48]) , (regs_regs_0_lpi_2[51:50]) , (regs_regs_0_lpi_2[53:52])
      , (regs_regs_0_lpi_2[55:54]) , (regs_regs_0_lpi_2[57:56]) , (regs_regs_0_lpi_2[59:58])
      , (regs_regs_0_lpi_2[61:60]) , (regs_regs_0_lpi_2[63:62]) , (regs_regs_0_lpi_2[65:64])
      , (regs_regs_0_lpi_2[67:66]) , (regs_regs_0_lpi_2[69:68]) , (regs_regs_0_lpi_2[71:70])
      , (regs_regs_0_lpi_2[73:72]) , (regs_regs_0_lpi_2[75:74]) , (regs_regs_0_lpi_2[77:76])
      , (regs_regs_0_lpi_2[79:78]) , (regs_regs_0_lpi_2[81:80]) , (regs_regs_0_lpi_2[83:82])
      , (regs_regs_0_lpi_2[85:84]) , (regs_regs_0_lpi_2[87:86]) , (regs_regs_0_lpi_2[89:88])
      , (regs_regs_0_lpi_2[91:90]) , (regs_regs_0_lpi_2[93:92]) , (regs_regs_0_lpi_2[95:94])
      , (regs_regs_0_lpi_2[97:96]) , (regs_regs_0_lpi_2[99:98]) , (regs_regs_0_lpi_2[101:100])
      , (regs_regs_0_lpi_2[103:102]) , (regs_regs_0_lpi_2[105:104]) , (regs_regs_0_lpi_2[107:106])
      , (regs_regs_0_lpi_2[109:108]) , (regs_regs_0_lpi_2[111:110]) , (regs_regs_0_lpi_2[113:112])
      , (regs_regs_0_lpi_2[115:114]) , (regs_regs_0_lpi_2[117:116]) , (regs_regs_0_lpi_2[119:118])
      , (regs_regs_0_lpi_2[121:120]) , (regs_regs_0_lpi_2[123:122]) , (regs_regs_0_lpi_2[125:124])
      , (regs_regs_0_lpi_2[127:126]) , (regs_regs_0_lpi_2[129:128]) , (regs_regs_0_lpi_2[131:130])
      , (regs_regs_0_lpi_2[133:132]) , (regs_regs_0_lpi_2[135:134]) , (regs_regs_0_lpi_2[137:136])
      , (regs_regs_0_lpi_2[139:138]) , (regs_regs_0_lpi_2[141:140]) , (regs_regs_0_lpi_2[143:142])
      , (regs_regs_0_lpi_2[145:144]) , (regs_regs_0_lpi_2[147:146]) , (regs_regs_0_lpi_2[149:148])
      , (regs_regs_1_lpi_2[1:0]) , (regs_regs_1_lpi_2[3:2]) , (regs_regs_1_lpi_2[5:4])
      , (regs_regs_1_lpi_2[7:6]) , (regs_regs_1_lpi_2[9:8]) , (regs_regs_1_lpi_2[11:10])
      , (regs_regs_1_lpi_2[13:12]) , (regs_regs_1_lpi_2[15:14]) , (regs_regs_1_lpi_2[17:16])
      , (regs_regs_1_lpi_2[19:18]) , (regs_regs_1_lpi_2[21:20]) , (regs_regs_1_lpi_2[23:22])
      , (regs_regs_1_lpi_2[25:24]) , (regs_regs_1_lpi_2[27:26]) , (regs_regs_1_lpi_2[29:28])
      , (regs_regs_1_lpi_2[31:30]) , (regs_regs_1_lpi_2[33:32]) , (regs_regs_1_lpi_2[35:34])
      , (regs_regs_1_lpi_2[37:36]) , (regs_regs_1_lpi_2[39:38]) , (regs_regs_1_lpi_2[41:40])
      , (regs_regs_1_lpi_2[43:42]) , (regs_regs_1_lpi_2[45:44]) , (regs_regs_1_lpi_2[47:46])
      , (regs_regs_1_lpi_2[49:48]) , (regs_regs_1_lpi_2[51:50]) , (regs_regs_1_lpi_2[53:52])
      , (regs_regs_1_lpi_2[55:54]) , (regs_regs_1_lpi_2[57:56]) , (regs_regs_1_lpi_2[59:58])
      , (regs_regs_1_lpi_2[61:60]) , (regs_regs_1_lpi_2[63:62]) , (regs_regs_1_lpi_2[65:64])
      , (regs_regs_1_lpi_2[67:66]) , (regs_regs_1_lpi_2[69:68]) , (regs_regs_1_lpi_2[71:70])
      , (regs_regs_1_lpi_2[73:72]) , (regs_regs_1_lpi_2[75:74]) , (regs_regs_1_lpi_2[77:76])
      , (regs_regs_1_lpi_2[79:78]) , (regs_regs_1_lpi_2[81:80]) , (regs_regs_1_lpi_2[83:82])
      , (regs_regs_1_lpi_2[85:84]) , (regs_regs_1_lpi_2[87:86]) , (regs_regs_1_lpi_2[89:88])
      , (regs_regs_1_lpi_2[91:90]) , (regs_regs_1_lpi_2[93:92]) , (regs_regs_1_lpi_2[95:94])
      , (regs_regs_1_lpi_2[97:96]) , (regs_regs_1_lpi_2[99:98]) , (regs_regs_1_lpi_2[101:100])
      , (regs_regs_1_lpi_2[103:102]) , (regs_regs_1_lpi_2[105:104]) , (regs_regs_1_lpi_2[107:106])
      , (regs_regs_1_lpi_2[109:108]) , (regs_regs_1_lpi_2[111:110]) , (regs_regs_1_lpi_2[113:112])
      , (regs_regs_1_lpi_2[115:114]) , (regs_regs_1_lpi_2[117:116]) , (regs_regs_1_lpi_2[119:118])
      , (regs_regs_1_lpi_2[121:120]) , (regs_regs_1_lpi_2[123:122]) , (regs_regs_1_lpi_2[125:124])
      , (regs_regs_1_lpi_2[127:126]) , (regs_regs_1_lpi_2[129:128]) , (regs_regs_1_lpi_2[131:130])
      , (regs_regs_1_lpi_2[133:132]) , (regs_regs_1_lpi_2[135:134]) , (regs_regs_1_lpi_2[137:136])
      , (regs_regs_1_lpi_2[139:138]) , (regs_regs_1_lpi_2[141:140]) , (regs_regs_1_lpi_2[143:142])
      , (regs_regs_1_lpi_2[145:144]) , (regs_regs_1_lpi_2[147:146]) , (regs_regs_1_lpi_2[149:148])
      , (regs_regs_2_lpi_2[1:0]) , (regs_regs_2_lpi_2[3:2]) , (regs_regs_2_lpi_2[5:4])
      , (regs_regs_2_lpi_2[7:6]) , (regs_regs_2_lpi_2[9:8]) , (regs_regs_2_lpi_2[11:10])
      , (regs_regs_2_lpi_2[13:12]) , (regs_regs_2_lpi_2[15:14]) , (regs_regs_2_lpi_2[17:16])
      , (regs_regs_2_lpi_2[19:18]) , (regs_regs_2_lpi_2[21:20]) , (regs_regs_2_lpi_2[23:22])
      , (regs_regs_2_lpi_2[25:24]) , (regs_regs_2_lpi_2[27:26]) , (regs_regs_2_lpi_2[29:28])
      , (regs_regs_2_lpi_2[31:30]) , (regs_regs_2_lpi_2[33:32]) , (regs_regs_2_lpi_2[35:34])
      , (regs_regs_2_lpi_2[37:36]) , (regs_regs_2_lpi_2[39:38]) , (regs_regs_2_lpi_2[41:40])
      , (regs_regs_2_lpi_2[43:42]) , (regs_regs_2_lpi_2[45:44]) , (regs_regs_2_lpi_2[47:46])
      , (regs_regs_2_lpi_2[49:48]) , (regs_regs_2_lpi_2[51:50]) , (regs_regs_2_lpi_2[53:52])
      , (regs_regs_2_lpi_2[55:54]) , (regs_regs_2_lpi_2[57:56]) , (regs_regs_2_lpi_2[59:58])
      , (regs_regs_2_lpi_2[61:60]) , (regs_regs_2_lpi_2[63:62]) , (regs_regs_2_lpi_2[65:64])
      , (regs_regs_2_lpi_2[67:66]) , (regs_regs_2_lpi_2[69:68]) , (regs_regs_2_lpi_2[71:70])
      , (regs_regs_2_lpi_2[73:72]) , (regs_regs_2_lpi_2[75:74]) , (regs_regs_2_lpi_2[77:76])
      , (regs_regs_2_lpi_2[79:78]) , (regs_regs_2_lpi_2[81:80]) , (regs_regs_2_lpi_2[83:82])
      , (regs_regs_2_lpi_2[85:84]) , (regs_regs_2_lpi_2[87:86]) , (regs_regs_2_lpi_2[89:88])
      , (regs_regs_2_lpi_2[91:90]) , (regs_regs_2_lpi_2[93:92]) , (regs_regs_2_lpi_2[95:94])
      , (regs_regs_2_lpi_2[97:96]) , (regs_regs_2_lpi_2[99:98]) , (regs_regs_2_lpi_2[101:100])
      , (regs_regs_2_lpi_2[103:102]) , (regs_regs_2_lpi_2[105:104]) , (regs_regs_2_lpi_2[107:106])
      , (regs_regs_2_lpi_2[109:108]) , (regs_regs_2_lpi_2[111:110]) , (regs_regs_2_lpi_2[113:112])
      , (regs_regs_2_lpi_2[115:114]) , (regs_regs_2_lpi_2[117:116]) , (regs_regs_2_lpi_2[119:118])
      , (regs_regs_2_lpi_2[121:120]) , (regs_regs_2_lpi_2[123:122]) , (regs_regs_2_lpi_2[125:124])
      , (regs_regs_2_lpi_2[127:126]) , (regs_regs_2_lpi_2[129:128]) , (regs_regs_2_lpi_2[131:130])
      , (regs_regs_2_lpi_2[133:132]) , (regs_regs_2_lpi_2[135:134]) , (regs_regs_2_lpi_2[137:136])
      , (regs_regs_2_lpi_2[139:138]) , (regs_regs_2_lpi_2[141:140]) , (regs_regs_2_lpi_2[143:142])
      , (regs_regs_2_lpi_2[145:144]) , (regs_regs_2_lpi_2[147:146]) , (regs_regs_2_lpi_2[149:148])
      , (regs_regs_3_lpi_2[1:0]) , (regs_regs_3_lpi_2[3:2]) , (regs_regs_3_lpi_2[5:4])
      , (regs_regs_3_lpi_2[7:6]) , (regs_regs_3_lpi_2[9:8]) , (regs_regs_3_lpi_2[11:10])
      , (regs_regs_3_lpi_2[13:12]) , (regs_regs_3_lpi_2[15:14]) , (regs_regs_3_lpi_2[17:16])
      , (regs_regs_3_lpi_2[19:18]) , (regs_regs_3_lpi_2[21:20]) , (regs_regs_3_lpi_2[23:22])
      , (regs_regs_3_lpi_2[25:24]) , (regs_regs_3_lpi_2[27:26]) , (regs_regs_3_lpi_2[29:28])
      , (regs_regs_3_lpi_2[31:30]) , (regs_regs_3_lpi_2[33:32]) , (regs_regs_3_lpi_2[35:34])
      , (regs_regs_3_lpi_2[37:36]) , (regs_regs_3_lpi_2[39:38]) , (regs_regs_3_lpi_2[41:40])
      , (regs_regs_3_lpi_2[43:42]) , (regs_regs_3_lpi_2[45:44]) , (regs_regs_3_lpi_2[47:46])
      , (regs_regs_3_lpi_2[49:48]) , (regs_regs_3_lpi_2[51:50]) , (regs_regs_3_lpi_2[53:52])
      , (regs_regs_3_lpi_2[55:54]) , (regs_regs_3_lpi_2[57:56]) , (regs_regs_3_lpi_2[59:58])
      , (regs_regs_3_lpi_2[61:60]) , (regs_regs_3_lpi_2[63:62]) , (regs_regs_3_lpi_2[65:64])
      , (regs_regs_3_lpi_2[67:66]) , (regs_regs_3_lpi_2[69:68]) , (regs_regs_3_lpi_2[71:70])
      , (regs_regs_3_lpi_2[73:72]) , (regs_regs_3_lpi_2[75:74]) , (regs_regs_3_lpi_2[77:76])
      , (regs_regs_3_lpi_2[79:78]) , (regs_regs_3_lpi_2[81:80]) , (regs_regs_3_lpi_2[83:82])
      , (regs_regs_3_lpi_2[85:84]) , (regs_regs_3_lpi_2[87:86]) , (regs_regs_3_lpi_2[89:88])
      , (regs_regs_3_lpi_2[91:90]) , (regs_regs_3_lpi_2[93:92]) , (regs_regs_3_lpi_2[95:94])
      , (regs_regs_3_lpi_2[97:96]) , (regs_regs_3_lpi_2[99:98]) , (regs_regs_3_lpi_2[101:100])
      , (regs_regs_3_lpi_2[103:102]) , (regs_regs_3_lpi_2[105:104]) , (regs_regs_3_lpi_2[107:106])
      , (regs_regs_3_lpi_2[109:108]) , (regs_regs_3_lpi_2[111:110]) , (regs_regs_3_lpi_2[113:112])
      , (regs_regs_3_lpi_2[115:114]) , (regs_regs_3_lpi_2[117:116]) , (regs_regs_3_lpi_2[119:118])
      , (regs_regs_3_lpi_2[121:120]) , (regs_regs_3_lpi_2[123:122]) , (regs_regs_3_lpi_2[125:124])
      , (regs_regs_3_lpi_2[127:126]) , (regs_regs_3_lpi_2[129:128]) , (regs_regs_3_lpi_2[131:130])
      , (regs_regs_3_lpi_2[133:132]) , (regs_regs_3_lpi_2[135:134]) , (regs_regs_3_lpi_2[137:136])
      , (regs_regs_3_lpi_2[139:138]) , (regs_regs_3_lpi_2[141:140]) , (regs_regs_3_lpi_2[143:142])
      , (regs_regs_3_lpi_2[145:144]) , (regs_regs_3_lpi_2[147:146]) , (regs_regs_3_lpi_2[149:148])
      , (regs_regs_4_lpi_2[1:0]) , (regs_regs_4_lpi_2[3:2]) , (regs_regs_4_lpi_2[5:4])
      , (regs_regs_4_lpi_2[7:6]) , (regs_regs_4_lpi_2[9:8]) , (regs_regs_4_lpi_2[11:10])
      , (regs_regs_4_lpi_2[13:12]) , (regs_regs_4_lpi_2[15:14]) , (regs_regs_4_lpi_2[17:16])
      , (regs_regs_4_lpi_2[19:18]) , (regs_regs_4_lpi_2[21:20]) , (regs_regs_4_lpi_2[23:22])
      , (regs_regs_4_lpi_2[25:24]) , (regs_regs_4_lpi_2[27:26]) , (regs_regs_4_lpi_2[29:28])
      , (regs_regs_4_lpi_2[31:30]) , (regs_regs_4_lpi_2[33:32]) , (regs_regs_4_lpi_2[35:34])
      , (regs_regs_4_lpi_2[37:36]) , (regs_regs_4_lpi_2[39:38]) , (regs_regs_4_lpi_2[41:40])
      , (regs_regs_4_lpi_2[43:42]) , (regs_regs_4_lpi_2[45:44]) , (regs_regs_4_lpi_2[47:46])
      , (regs_regs_4_lpi_2[49:48]) , (regs_regs_4_lpi_2[51:50]) , (regs_regs_4_lpi_2[53:52])
      , (regs_regs_4_lpi_2[55:54]) , (regs_regs_4_lpi_2[57:56]) , (regs_regs_4_lpi_2[59:58])
      , (regs_regs_4_lpi_2[61:60]) , (regs_regs_4_lpi_2[63:62]) , (regs_regs_4_lpi_2[65:64])
      , (regs_regs_4_lpi_2[67:66]) , (regs_regs_4_lpi_2[69:68]) , (regs_regs_4_lpi_2[71:70])
      , (regs_regs_4_lpi_2[73:72]) , (regs_regs_4_lpi_2[75:74]) , (regs_regs_4_lpi_2[77:76])
      , (regs_regs_4_lpi_2[79:78]) , (regs_regs_4_lpi_2[81:80]) , (regs_regs_4_lpi_2[83:82])
      , (regs_regs_4_lpi_2[85:84]) , (regs_regs_4_lpi_2[87:86]) , (regs_regs_4_lpi_2[89:88])
      , (regs_regs_4_lpi_2[91:90]) , (regs_regs_4_lpi_2[93:92]) , (regs_regs_4_lpi_2[95:94])
      , (regs_regs_4_lpi_2[97:96]) , (regs_regs_4_lpi_2[99:98]) , (regs_regs_4_lpi_2[101:100])
      , (regs_regs_4_lpi_2[103:102]) , (regs_regs_4_lpi_2[105:104]) , (regs_regs_4_lpi_2[107:106])
      , (regs_regs_4_lpi_2[109:108]) , (regs_regs_4_lpi_2[111:110]) , (regs_regs_4_lpi_2[113:112])
      , (regs_regs_4_lpi_2[115:114]) , (regs_regs_4_lpi_2[117:116]) , (regs_regs_4_lpi_2[119:118])
      , (regs_regs_4_lpi_2[121:120]) , (regs_regs_4_lpi_2[123:122]) , (regs_regs_4_lpi_2[125:124])
      , (regs_regs_4_lpi_2[127:126]) , (regs_regs_4_lpi_2[129:128]) , (regs_regs_4_lpi_2[131:130])
      , (regs_regs_4_lpi_2[133:132]) , (regs_regs_4_lpi_2[135:134]) , (regs_regs_4_lpi_2[137:136])
      , (regs_regs_4_lpi_2[139:138]) , (regs_regs_4_lpi_2[141:140]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg9 = MUX_v_2_512_2({(regs_regs_0_lpi_2[19:18]) , (regs_regs_0_lpi_2[21:20])
      , (regs_regs_0_lpi_2[23:22]) , (regs_regs_0_lpi_2[25:24]) , (regs_regs_0_lpi_2[27:26])
      , (regs_regs_0_lpi_2[29:28]) , (regs_regs_0_lpi_2[31:30]) , (regs_regs_0_lpi_2[33:32])
      , (regs_regs_0_lpi_2[35:34]) , (regs_regs_0_lpi_2[37:36]) , (regs_regs_0_lpi_2[39:38])
      , (regs_regs_0_lpi_2[41:40]) , (regs_regs_0_lpi_2[43:42]) , (regs_regs_0_lpi_2[45:44])
      , (regs_regs_0_lpi_2[47:46]) , (regs_regs_0_lpi_2[49:48]) , (regs_regs_0_lpi_2[51:50])
      , (regs_regs_0_lpi_2[53:52]) , (regs_regs_0_lpi_2[55:54]) , (regs_regs_0_lpi_2[57:56])
      , (regs_regs_0_lpi_2[59:58]) , (regs_regs_0_lpi_2[61:60]) , (regs_regs_0_lpi_2[63:62])
      , (regs_regs_0_lpi_2[65:64]) , (regs_regs_0_lpi_2[67:66]) , (regs_regs_0_lpi_2[69:68])
      , (regs_regs_0_lpi_2[71:70]) , (regs_regs_0_lpi_2[73:72]) , (regs_regs_0_lpi_2[75:74])
      , (regs_regs_0_lpi_2[77:76]) , (regs_regs_0_lpi_2[79:78]) , (regs_regs_0_lpi_2[81:80])
      , (regs_regs_0_lpi_2[83:82]) , (regs_regs_0_lpi_2[85:84]) , (regs_regs_0_lpi_2[87:86])
      , (regs_regs_0_lpi_2[89:88]) , (regs_regs_0_lpi_2[91:90]) , (regs_regs_0_lpi_2[93:92])
      , (regs_regs_0_lpi_2[95:94]) , (regs_regs_0_lpi_2[97:96]) , (regs_regs_0_lpi_2[99:98])
      , (regs_regs_0_lpi_2[101:100]) , (regs_regs_0_lpi_2[103:102]) , (regs_regs_0_lpi_2[105:104])
      , (regs_regs_0_lpi_2[107:106]) , (regs_regs_0_lpi_2[109:108]) , (regs_regs_0_lpi_2[111:110])
      , (regs_regs_0_lpi_2[113:112]) , (regs_regs_0_lpi_2[115:114]) , (regs_regs_0_lpi_2[117:116])
      , (regs_regs_0_lpi_2[119:118]) , (regs_regs_0_lpi_2[121:120]) , (regs_regs_0_lpi_2[123:122])
      , (regs_regs_0_lpi_2[125:124]) , (regs_regs_0_lpi_2[127:126]) , (regs_regs_0_lpi_2[129:128])
      , (regs_regs_0_lpi_2[131:130]) , (regs_regs_0_lpi_2[133:132]) , (regs_regs_0_lpi_2[135:134])
      , (regs_regs_0_lpi_2[137:136]) , (regs_regs_0_lpi_2[139:138]) , (regs_regs_0_lpi_2[141:140])
      , (regs_regs_0_lpi_2[143:142]) , (regs_regs_0_lpi_2[145:144]) , (regs_regs_0_lpi_2[147:146])
      , (regs_regs_0_lpi_2[149:148]) , (regs_regs_1_lpi_2[1:0]) , (regs_regs_1_lpi_2[3:2])
      , (regs_regs_1_lpi_2[5:4]) , (regs_regs_1_lpi_2[7:6]) , (regs_regs_1_lpi_2[9:8])
      , (regs_regs_1_lpi_2[11:10]) , (regs_regs_1_lpi_2[13:12]) , (regs_regs_1_lpi_2[15:14])
      , (regs_regs_1_lpi_2[17:16]) , (regs_regs_1_lpi_2[19:18]) , (regs_regs_1_lpi_2[21:20])
      , (regs_regs_1_lpi_2[23:22]) , (regs_regs_1_lpi_2[25:24]) , (regs_regs_1_lpi_2[27:26])
      , (regs_regs_1_lpi_2[29:28]) , (regs_regs_1_lpi_2[31:30]) , (regs_regs_1_lpi_2[33:32])
      , (regs_regs_1_lpi_2[35:34]) , (regs_regs_1_lpi_2[37:36]) , (regs_regs_1_lpi_2[39:38])
      , (regs_regs_1_lpi_2[41:40]) , (regs_regs_1_lpi_2[43:42]) , (regs_regs_1_lpi_2[45:44])
      , (regs_regs_1_lpi_2[47:46]) , (regs_regs_1_lpi_2[49:48]) , (regs_regs_1_lpi_2[51:50])
      , (regs_regs_1_lpi_2[53:52]) , (regs_regs_1_lpi_2[55:54]) , (regs_regs_1_lpi_2[57:56])
      , (regs_regs_1_lpi_2[59:58]) , (regs_regs_1_lpi_2[61:60]) , (regs_regs_1_lpi_2[63:62])
      , (regs_regs_1_lpi_2[65:64]) , (regs_regs_1_lpi_2[67:66]) , (regs_regs_1_lpi_2[69:68])
      , (regs_regs_1_lpi_2[71:70]) , (regs_regs_1_lpi_2[73:72]) , (regs_regs_1_lpi_2[75:74])
      , (regs_regs_1_lpi_2[77:76]) , (regs_regs_1_lpi_2[79:78]) , (regs_regs_1_lpi_2[81:80])
      , (regs_regs_1_lpi_2[83:82]) , (regs_regs_1_lpi_2[85:84]) , (regs_regs_1_lpi_2[87:86])
      , (regs_regs_1_lpi_2[89:88]) , (regs_regs_1_lpi_2[91:90]) , (regs_regs_1_lpi_2[93:92])
      , (regs_regs_1_lpi_2[95:94]) , (regs_regs_1_lpi_2[97:96]) , (regs_regs_1_lpi_2[99:98])
      , (regs_regs_1_lpi_2[101:100]) , (regs_regs_1_lpi_2[103:102]) , (regs_regs_1_lpi_2[105:104])
      , (regs_regs_1_lpi_2[107:106]) , (regs_regs_1_lpi_2[109:108]) , (regs_regs_1_lpi_2[111:110])
      , (regs_regs_1_lpi_2[113:112]) , (regs_regs_1_lpi_2[115:114]) , (regs_regs_1_lpi_2[117:116])
      , (regs_regs_1_lpi_2[119:118]) , (regs_regs_1_lpi_2[121:120]) , (regs_regs_1_lpi_2[123:122])
      , (regs_regs_1_lpi_2[125:124]) , (regs_regs_1_lpi_2[127:126]) , (regs_regs_1_lpi_2[129:128])
      , (regs_regs_1_lpi_2[131:130]) , (regs_regs_1_lpi_2[133:132]) , (regs_regs_1_lpi_2[135:134])
      , (regs_regs_1_lpi_2[137:136]) , (regs_regs_1_lpi_2[139:138]) , (regs_regs_1_lpi_2[141:140])
      , (regs_regs_1_lpi_2[143:142]) , (regs_regs_1_lpi_2[145:144]) , (regs_regs_1_lpi_2[147:146])
      , (regs_regs_1_lpi_2[149:148]) , (regs_regs_2_lpi_2[1:0]) , (regs_regs_2_lpi_2[3:2])
      , (regs_regs_2_lpi_2[5:4]) , (regs_regs_2_lpi_2[7:6]) , (regs_regs_2_lpi_2[9:8])
      , (regs_regs_2_lpi_2[11:10]) , (regs_regs_2_lpi_2[13:12]) , (regs_regs_2_lpi_2[15:14])
      , (regs_regs_2_lpi_2[17:16]) , (regs_regs_2_lpi_2[19:18]) , (regs_regs_2_lpi_2[21:20])
      , (regs_regs_2_lpi_2[23:22]) , (regs_regs_2_lpi_2[25:24]) , (regs_regs_2_lpi_2[27:26])
      , (regs_regs_2_lpi_2[29:28]) , (regs_regs_2_lpi_2[31:30]) , (regs_regs_2_lpi_2[33:32])
      , (regs_regs_2_lpi_2[35:34]) , (regs_regs_2_lpi_2[37:36]) , (regs_regs_2_lpi_2[39:38])
      , (regs_regs_2_lpi_2[41:40]) , (regs_regs_2_lpi_2[43:42]) , (regs_regs_2_lpi_2[45:44])
      , (regs_regs_2_lpi_2[47:46]) , (regs_regs_2_lpi_2[49:48]) , (regs_regs_2_lpi_2[51:50])
      , (regs_regs_2_lpi_2[53:52]) , (regs_regs_2_lpi_2[55:54]) , (regs_regs_2_lpi_2[57:56])
      , (regs_regs_2_lpi_2[59:58]) , (regs_regs_2_lpi_2[61:60]) , (regs_regs_2_lpi_2[63:62])
      , (regs_regs_2_lpi_2[65:64]) , (regs_regs_2_lpi_2[67:66]) , (regs_regs_2_lpi_2[69:68])
      , (regs_regs_2_lpi_2[71:70]) , (regs_regs_2_lpi_2[73:72]) , (regs_regs_2_lpi_2[75:74])
      , (regs_regs_2_lpi_2[77:76]) , (regs_regs_2_lpi_2[79:78]) , (regs_regs_2_lpi_2[81:80])
      , (regs_regs_2_lpi_2[83:82]) , (regs_regs_2_lpi_2[85:84]) , (regs_regs_2_lpi_2[87:86])
      , (regs_regs_2_lpi_2[89:88]) , (regs_regs_2_lpi_2[91:90]) , (regs_regs_2_lpi_2[93:92])
      , (regs_regs_2_lpi_2[95:94]) , (regs_regs_2_lpi_2[97:96]) , (regs_regs_2_lpi_2[99:98])
      , (regs_regs_2_lpi_2[101:100]) , (regs_regs_2_lpi_2[103:102]) , (regs_regs_2_lpi_2[105:104])
      , (regs_regs_2_lpi_2[107:106]) , (regs_regs_2_lpi_2[109:108]) , (regs_regs_2_lpi_2[111:110])
      , (regs_regs_2_lpi_2[113:112]) , (regs_regs_2_lpi_2[115:114]) , (regs_regs_2_lpi_2[117:116])
      , (regs_regs_2_lpi_2[119:118]) , (regs_regs_2_lpi_2[121:120]) , (regs_regs_2_lpi_2[123:122])
      , (regs_regs_2_lpi_2[125:124]) , (regs_regs_2_lpi_2[127:126]) , (regs_regs_2_lpi_2[129:128])
      , (regs_regs_2_lpi_2[131:130]) , (regs_regs_2_lpi_2[133:132]) , (regs_regs_2_lpi_2[135:134])
      , (regs_regs_2_lpi_2[137:136]) , (regs_regs_2_lpi_2[139:138]) , (regs_regs_2_lpi_2[141:140])
      , (regs_regs_2_lpi_2[143:142]) , (regs_regs_2_lpi_2[145:144]) , (regs_regs_2_lpi_2[147:146])
      , (regs_regs_2_lpi_2[149:148]) , (regs_regs_3_lpi_2[1:0]) , (regs_regs_3_lpi_2[3:2])
      , (regs_regs_3_lpi_2[5:4]) , (regs_regs_3_lpi_2[7:6]) , (regs_regs_3_lpi_2[9:8])
      , (regs_regs_3_lpi_2[11:10]) , (regs_regs_3_lpi_2[13:12]) , (regs_regs_3_lpi_2[15:14])
      , (regs_regs_3_lpi_2[17:16]) , (regs_regs_3_lpi_2[19:18]) , (regs_regs_3_lpi_2[21:20])
      , (regs_regs_3_lpi_2[23:22]) , (regs_regs_3_lpi_2[25:24]) , (regs_regs_3_lpi_2[27:26])
      , (regs_regs_3_lpi_2[29:28]) , (regs_regs_3_lpi_2[31:30]) , (regs_regs_3_lpi_2[33:32])
      , (regs_regs_3_lpi_2[35:34]) , (regs_regs_3_lpi_2[37:36]) , (regs_regs_3_lpi_2[39:38])
      , (regs_regs_3_lpi_2[41:40]) , (regs_regs_3_lpi_2[43:42]) , (regs_regs_3_lpi_2[45:44])
      , (regs_regs_3_lpi_2[47:46]) , (regs_regs_3_lpi_2[49:48]) , (regs_regs_3_lpi_2[51:50])
      , (regs_regs_3_lpi_2[53:52]) , (regs_regs_3_lpi_2[55:54]) , (regs_regs_3_lpi_2[57:56])
      , (regs_regs_3_lpi_2[59:58]) , (regs_regs_3_lpi_2[61:60]) , (regs_regs_3_lpi_2[63:62])
      , (regs_regs_3_lpi_2[65:64]) , (regs_regs_3_lpi_2[67:66]) , (regs_regs_3_lpi_2[69:68])
      , (regs_regs_3_lpi_2[71:70]) , (regs_regs_3_lpi_2[73:72]) , (regs_regs_3_lpi_2[75:74])
      , (regs_regs_3_lpi_2[77:76]) , (regs_regs_3_lpi_2[79:78]) , (regs_regs_3_lpi_2[81:80])
      , (regs_regs_3_lpi_2[83:82]) , (regs_regs_3_lpi_2[85:84]) , (regs_regs_3_lpi_2[87:86])
      , (regs_regs_3_lpi_2[89:88]) , (regs_regs_3_lpi_2[91:90]) , (regs_regs_3_lpi_2[93:92])
      , (regs_regs_3_lpi_2[95:94]) , (regs_regs_3_lpi_2[97:96]) , (regs_regs_3_lpi_2[99:98])
      , (regs_regs_3_lpi_2[101:100]) , (regs_regs_3_lpi_2[103:102]) , (regs_regs_3_lpi_2[105:104])
      , (regs_regs_3_lpi_2[107:106]) , (regs_regs_3_lpi_2[109:108]) , (regs_regs_3_lpi_2[111:110])
      , (regs_regs_3_lpi_2[113:112]) , (regs_regs_3_lpi_2[115:114]) , (regs_regs_3_lpi_2[117:116])
      , (regs_regs_3_lpi_2[119:118]) , (regs_regs_3_lpi_2[121:120]) , (regs_regs_3_lpi_2[123:122])
      , (regs_regs_3_lpi_2[125:124]) , (regs_regs_3_lpi_2[127:126]) , (regs_regs_3_lpi_2[129:128])
      , (regs_regs_3_lpi_2[131:130]) , (regs_regs_3_lpi_2[133:132]) , (regs_regs_3_lpi_2[135:134])
      , (regs_regs_3_lpi_2[137:136]) , (regs_regs_3_lpi_2[139:138]) , (regs_regs_3_lpi_2[141:140])
      , (regs_regs_3_lpi_2[143:142]) , (regs_regs_3_lpi_2[145:144]) , (regs_regs_3_lpi_2[147:146])
      , (regs_regs_3_lpi_2[149:148]) , (regs_regs_4_lpi_2[1:0]) , (regs_regs_4_lpi_2[3:2])
      , (regs_regs_4_lpi_2[5:4]) , (regs_regs_4_lpi_2[7:6]) , (regs_regs_4_lpi_2[9:8])
      , (regs_regs_4_lpi_2[11:10]) , (regs_regs_4_lpi_2[13:12]) , (regs_regs_4_lpi_2[15:14])
      , (regs_regs_4_lpi_2[17:16]) , (regs_regs_4_lpi_2[19:18]) , (regs_regs_4_lpi_2[21:20])
      , (regs_regs_4_lpi_2[23:22]) , (regs_regs_4_lpi_2[25:24]) , (regs_regs_4_lpi_2[27:26])
      , (regs_regs_4_lpi_2[29:28]) , (regs_regs_4_lpi_2[31:30]) , (regs_regs_4_lpi_2[33:32])
      , (regs_regs_4_lpi_2[35:34]) , (regs_regs_4_lpi_2[37:36]) , (regs_regs_4_lpi_2[39:38])
      , (regs_regs_4_lpi_2[41:40]) , (regs_regs_4_lpi_2[43:42]) , (regs_regs_4_lpi_2[45:44])
      , (regs_regs_4_lpi_2[47:46]) , (regs_regs_4_lpi_2[49:48]) , (regs_regs_4_lpi_2[51:50])
      , (regs_regs_4_lpi_2[53:52]) , (regs_regs_4_lpi_2[55:54]) , (regs_regs_4_lpi_2[57:56])
      , (regs_regs_4_lpi_2[59:58]) , (regs_regs_4_lpi_2[61:60]) , (regs_regs_4_lpi_2[63:62])
      , (regs_regs_4_lpi_2[65:64]) , (regs_regs_4_lpi_2[67:66]) , (regs_regs_4_lpi_2[69:68])
      , (regs_regs_4_lpi_2[71:70]) , (regs_regs_4_lpi_2[73:72]) , (regs_regs_4_lpi_2[75:74])
      , (regs_regs_4_lpi_2[77:76]) , (regs_regs_4_lpi_2[79:78]) , (regs_regs_4_lpi_2[81:80])
      , (regs_regs_4_lpi_2[83:82]) , (regs_regs_4_lpi_2[85:84]) , (regs_regs_4_lpi_2[87:86])
      , (regs_regs_4_lpi_2[89:88]) , (regs_regs_4_lpi_2[91:90]) , (regs_regs_4_lpi_2[93:92])
      , (regs_regs_4_lpi_2[95:94]) , (regs_regs_4_lpi_2[97:96]) , (regs_regs_4_lpi_2[99:98])
      , (regs_regs_4_lpi_2[101:100]) , (regs_regs_4_lpi_2[103:102]) , (regs_regs_4_lpi_2[105:104])
      , (regs_regs_4_lpi_2[107:106]) , (regs_regs_4_lpi_2[109:108]) , (regs_regs_4_lpi_2[111:110])
      , (regs_regs_4_lpi_2[113:112]) , (regs_regs_4_lpi_2[115:114]) , (regs_regs_4_lpi_2[117:116])
      , (regs_regs_4_lpi_2[119:118]) , (regs_regs_4_lpi_2[121:120]) , (regs_regs_4_lpi_2[123:122])
      , (regs_regs_4_lpi_2[125:124]) , (regs_regs_4_lpi_2[127:126]) , (regs_regs_4_lpi_2[129:128])
      , (regs_regs_4_lpi_2[131:130]) , (regs_regs_4_lpi_2[133:132]) , (regs_regs_4_lpi_2[135:134])
      , (regs_regs_4_lpi_2[137:136]) , (regs_regs_4_lpi_2[139:138]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg8 = MUX_v_2_512_2({(regs_regs_0_lpi_2[17:16]) , (regs_regs_0_lpi_2[19:18])
      , (regs_regs_0_lpi_2[21:20]) , (regs_regs_0_lpi_2[23:22]) , (regs_regs_0_lpi_2[25:24])
      , (regs_regs_0_lpi_2[27:26]) , (regs_regs_0_lpi_2[29:28]) , (regs_regs_0_lpi_2[31:30])
      , (regs_regs_0_lpi_2[33:32]) , (regs_regs_0_lpi_2[35:34]) , (regs_regs_0_lpi_2[37:36])
      , (regs_regs_0_lpi_2[39:38]) , (regs_regs_0_lpi_2[41:40]) , (regs_regs_0_lpi_2[43:42])
      , (regs_regs_0_lpi_2[45:44]) , (regs_regs_0_lpi_2[47:46]) , (regs_regs_0_lpi_2[49:48])
      , (regs_regs_0_lpi_2[51:50]) , (regs_regs_0_lpi_2[53:52]) , (regs_regs_0_lpi_2[55:54])
      , (regs_regs_0_lpi_2[57:56]) , (regs_regs_0_lpi_2[59:58]) , (regs_regs_0_lpi_2[61:60])
      , (regs_regs_0_lpi_2[63:62]) , (regs_regs_0_lpi_2[65:64]) , (regs_regs_0_lpi_2[67:66])
      , (regs_regs_0_lpi_2[69:68]) , (regs_regs_0_lpi_2[71:70]) , (regs_regs_0_lpi_2[73:72])
      , (regs_regs_0_lpi_2[75:74]) , (regs_regs_0_lpi_2[77:76]) , (regs_regs_0_lpi_2[79:78])
      , (regs_regs_0_lpi_2[81:80]) , (regs_regs_0_lpi_2[83:82]) , (regs_regs_0_lpi_2[85:84])
      , (regs_regs_0_lpi_2[87:86]) , (regs_regs_0_lpi_2[89:88]) , (regs_regs_0_lpi_2[91:90])
      , (regs_regs_0_lpi_2[93:92]) , (regs_regs_0_lpi_2[95:94]) , (regs_regs_0_lpi_2[97:96])
      , (regs_regs_0_lpi_2[99:98]) , (regs_regs_0_lpi_2[101:100]) , (regs_regs_0_lpi_2[103:102])
      , (regs_regs_0_lpi_2[105:104]) , (regs_regs_0_lpi_2[107:106]) , (regs_regs_0_lpi_2[109:108])
      , (regs_regs_0_lpi_2[111:110]) , (regs_regs_0_lpi_2[113:112]) , (regs_regs_0_lpi_2[115:114])
      , (regs_regs_0_lpi_2[117:116]) , (regs_regs_0_lpi_2[119:118]) , (regs_regs_0_lpi_2[121:120])
      , (regs_regs_0_lpi_2[123:122]) , (regs_regs_0_lpi_2[125:124]) , (regs_regs_0_lpi_2[127:126])
      , (regs_regs_0_lpi_2[129:128]) , (regs_regs_0_lpi_2[131:130]) , (regs_regs_0_lpi_2[133:132])
      , (regs_regs_0_lpi_2[135:134]) , (regs_regs_0_lpi_2[137:136]) , (regs_regs_0_lpi_2[139:138])
      , (regs_regs_0_lpi_2[141:140]) , (regs_regs_0_lpi_2[143:142]) , (regs_regs_0_lpi_2[145:144])
      , (regs_regs_0_lpi_2[147:146]) , (regs_regs_0_lpi_2[149:148]) , (regs_regs_1_lpi_2[1:0])
      , (regs_regs_1_lpi_2[3:2]) , (regs_regs_1_lpi_2[5:4]) , (regs_regs_1_lpi_2[7:6])
      , (regs_regs_1_lpi_2[9:8]) , (regs_regs_1_lpi_2[11:10]) , (regs_regs_1_lpi_2[13:12])
      , (regs_regs_1_lpi_2[15:14]) , (regs_regs_1_lpi_2[17:16]) , (regs_regs_1_lpi_2[19:18])
      , (regs_regs_1_lpi_2[21:20]) , (regs_regs_1_lpi_2[23:22]) , (regs_regs_1_lpi_2[25:24])
      , (regs_regs_1_lpi_2[27:26]) , (regs_regs_1_lpi_2[29:28]) , (regs_regs_1_lpi_2[31:30])
      , (regs_regs_1_lpi_2[33:32]) , (regs_regs_1_lpi_2[35:34]) , (regs_regs_1_lpi_2[37:36])
      , (regs_regs_1_lpi_2[39:38]) , (regs_regs_1_lpi_2[41:40]) , (regs_regs_1_lpi_2[43:42])
      , (regs_regs_1_lpi_2[45:44]) , (regs_regs_1_lpi_2[47:46]) , (regs_regs_1_lpi_2[49:48])
      , (regs_regs_1_lpi_2[51:50]) , (regs_regs_1_lpi_2[53:52]) , (regs_regs_1_lpi_2[55:54])
      , (regs_regs_1_lpi_2[57:56]) , (regs_regs_1_lpi_2[59:58]) , (regs_regs_1_lpi_2[61:60])
      , (regs_regs_1_lpi_2[63:62]) , (regs_regs_1_lpi_2[65:64]) , (regs_regs_1_lpi_2[67:66])
      , (regs_regs_1_lpi_2[69:68]) , (regs_regs_1_lpi_2[71:70]) , (regs_regs_1_lpi_2[73:72])
      , (regs_regs_1_lpi_2[75:74]) , (regs_regs_1_lpi_2[77:76]) , (regs_regs_1_lpi_2[79:78])
      , (regs_regs_1_lpi_2[81:80]) , (regs_regs_1_lpi_2[83:82]) , (regs_regs_1_lpi_2[85:84])
      , (regs_regs_1_lpi_2[87:86]) , (regs_regs_1_lpi_2[89:88]) , (regs_regs_1_lpi_2[91:90])
      , (regs_regs_1_lpi_2[93:92]) , (regs_regs_1_lpi_2[95:94]) , (regs_regs_1_lpi_2[97:96])
      , (regs_regs_1_lpi_2[99:98]) , (regs_regs_1_lpi_2[101:100]) , (regs_regs_1_lpi_2[103:102])
      , (regs_regs_1_lpi_2[105:104]) , (regs_regs_1_lpi_2[107:106]) , (regs_regs_1_lpi_2[109:108])
      , (regs_regs_1_lpi_2[111:110]) , (regs_regs_1_lpi_2[113:112]) , (regs_regs_1_lpi_2[115:114])
      , (regs_regs_1_lpi_2[117:116]) , (regs_regs_1_lpi_2[119:118]) , (regs_regs_1_lpi_2[121:120])
      , (regs_regs_1_lpi_2[123:122]) , (regs_regs_1_lpi_2[125:124]) , (regs_regs_1_lpi_2[127:126])
      , (regs_regs_1_lpi_2[129:128]) , (regs_regs_1_lpi_2[131:130]) , (regs_regs_1_lpi_2[133:132])
      , (regs_regs_1_lpi_2[135:134]) , (regs_regs_1_lpi_2[137:136]) , (regs_regs_1_lpi_2[139:138])
      , (regs_regs_1_lpi_2[141:140]) , (regs_regs_1_lpi_2[143:142]) , (regs_regs_1_lpi_2[145:144])
      , (regs_regs_1_lpi_2[147:146]) , (regs_regs_1_lpi_2[149:148]) , (regs_regs_2_lpi_2[1:0])
      , (regs_regs_2_lpi_2[3:2]) , (regs_regs_2_lpi_2[5:4]) , (regs_regs_2_lpi_2[7:6])
      , (regs_regs_2_lpi_2[9:8]) , (regs_regs_2_lpi_2[11:10]) , (regs_regs_2_lpi_2[13:12])
      , (regs_regs_2_lpi_2[15:14]) , (regs_regs_2_lpi_2[17:16]) , (regs_regs_2_lpi_2[19:18])
      , (regs_regs_2_lpi_2[21:20]) , (regs_regs_2_lpi_2[23:22]) , (regs_regs_2_lpi_2[25:24])
      , (regs_regs_2_lpi_2[27:26]) , (regs_regs_2_lpi_2[29:28]) , (regs_regs_2_lpi_2[31:30])
      , (regs_regs_2_lpi_2[33:32]) , (regs_regs_2_lpi_2[35:34]) , (regs_regs_2_lpi_2[37:36])
      , (regs_regs_2_lpi_2[39:38]) , (regs_regs_2_lpi_2[41:40]) , (regs_regs_2_lpi_2[43:42])
      , (regs_regs_2_lpi_2[45:44]) , (regs_regs_2_lpi_2[47:46]) , (regs_regs_2_lpi_2[49:48])
      , (regs_regs_2_lpi_2[51:50]) , (regs_regs_2_lpi_2[53:52]) , (regs_regs_2_lpi_2[55:54])
      , (regs_regs_2_lpi_2[57:56]) , (regs_regs_2_lpi_2[59:58]) , (regs_regs_2_lpi_2[61:60])
      , (regs_regs_2_lpi_2[63:62]) , (regs_regs_2_lpi_2[65:64]) , (regs_regs_2_lpi_2[67:66])
      , (regs_regs_2_lpi_2[69:68]) , (regs_regs_2_lpi_2[71:70]) , (regs_regs_2_lpi_2[73:72])
      , (regs_regs_2_lpi_2[75:74]) , (regs_regs_2_lpi_2[77:76]) , (regs_regs_2_lpi_2[79:78])
      , (regs_regs_2_lpi_2[81:80]) , (regs_regs_2_lpi_2[83:82]) , (regs_regs_2_lpi_2[85:84])
      , (regs_regs_2_lpi_2[87:86]) , (regs_regs_2_lpi_2[89:88]) , (regs_regs_2_lpi_2[91:90])
      , (regs_regs_2_lpi_2[93:92]) , (regs_regs_2_lpi_2[95:94]) , (regs_regs_2_lpi_2[97:96])
      , (regs_regs_2_lpi_2[99:98]) , (regs_regs_2_lpi_2[101:100]) , (regs_regs_2_lpi_2[103:102])
      , (regs_regs_2_lpi_2[105:104]) , (regs_regs_2_lpi_2[107:106]) , (regs_regs_2_lpi_2[109:108])
      , (regs_regs_2_lpi_2[111:110]) , (regs_regs_2_lpi_2[113:112]) , (regs_regs_2_lpi_2[115:114])
      , (regs_regs_2_lpi_2[117:116]) , (regs_regs_2_lpi_2[119:118]) , (regs_regs_2_lpi_2[121:120])
      , (regs_regs_2_lpi_2[123:122]) , (regs_regs_2_lpi_2[125:124]) , (regs_regs_2_lpi_2[127:126])
      , (regs_regs_2_lpi_2[129:128]) , (regs_regs_2_lpi_2[131:130]) , (regs_regs_2_lpi_2[133:132])
      , (regs_regs_2_lpi_2[135:134]) , (regs_regs_2_lpi_2[137:136]) , (regs_regs_2_lpi_2[139:138])
      , (regs_regs_2_lpi_2[141:140]) , (regs_regs_2_lpi_2[143:142]) , (regs_regs_2_lpi_2[145:144])
      , (regs_regs_2_lpi_2[147:146]) , (regs_regs_2_lpi_2[149:148]) , (regs_regs_3_lpi_2[1:0])
      , (regs_regs_3_lpi_2[3:2]) , (regs_regs_3_lpi_2[5:4]) , (regs_regs_3_lpi_2[7:6])
      , (regs_regs_3_lpi_2[9:8]) , (regs_regs_3_lpi_2[11:10]) , (regs_regs_3_lpi_2[13:12])
      , (regs_regs_3_lpi_2[15:14]) , (regs_regs_3_lpi_2[17:16]) , (regs_regs_3_lpi_2[19:18])
      , (regs_regs_3_lpi_2[21:20]) , (regs_regs_3_lpi_2[23:22]) , (regs_regs_3_lpi_2[25:24])
      , (regs_regs_3_lpi_2[27:26]) , (regs_regs_3_lpi_2[29:28]) , (regs_regs_3_lpi_2[31:30])
      , (regs_regs_3_lpi_2[33:32]) , (regs_regs_3_lpi_2[35:34]) , (regs_regs_3_lpi_2[37:36])
      , (regs_regs_3_lpi_2[39:38]) , (regs_regs_3_lpi_2[41:40]) , (regs_regs_3_lpi_2[43:42])
      , (regs_regs_3_lpi_2[45:44]) , (regs_regs_3_lpi_2[47:46]) , (regs_regs_3_lpi_2[49:48])
      , (regs_regs_3_lpi_2[51:50]) , (regs_regs_3_lpi_2[53:52]) , (regs_regs_3_lpi_2[55:54])
      , (regs_regs_3_lpi_2[57:56]) , (regs_regs_3_lpi_2[59:58]) , (regs_regs_3_lpi_2[61:60])
      , (regs_regs_3_lpi_2[63:62]) , (regs_regs_3_lpi_2[65:64]) , (regs_regs_3_lpi_2[67:66])
      , (regs_regs_3_lpi_2[69:68]) , (regs_regs_3_lpi_2[71:70]) , (regs_regs_3_lpi_2[73:72])
      , (regs_regs_3_lpi_2[75:74]) , (regs_regs_3_lpi_2[77:76]) , (regs_regs_3_lpi_2[79:78])
      , (regs_regs_3_lpi_2[81:80]) , (regs_regs_3_lpi_2[83:82]) , (regs_regs_3_lpi_2[85:84])
      , (regs_regs_3_lpi_2[87:86]) , (regs_regs_3_lpi_2[89:88]) , (regs_regs_3_lpi_2[91:90])
      , (regs_regs_3_lpi_2[93:92]) , (regs_regs_3_lpi_2[95:94]) , (regs_regs_3_lpi_2[97:96])
      , (regs_regs_3_lpi_2[99:98]) , (regs_regs_3_lpi_2[101:100]) , (regs_regs_3_lpi_2[103:102])
      , (regs_regs_3_lpi_2[105:104]) , (regs_regs_3_lpi_2[107:106]) , (regs_regs_3_lpi_2[109:108])
      , (regs_regs_3_lpi_2[111:110]) , (regs_regs_3_lpi_2[113:112]) , (regs_regs_3_lpi_2[115:114])
      , (regs_regs_3_lpi_2[117:116]) , (regs_regs_3_lpi_2[119:118]) , (regs_regs_3_lpi_2[121:120])
      , (regs_regs_3_lpi_2[123:122]) , (regs_regs_3_lpi_2[125:124]) , (regs_regs_3_lpi_2[127:126])
      , (regs_regs_3_lpi_2[129:128]) , (regs_regs_3_lpi_2[131:130]) , (regs_regs_3_lpi_2[133:132])
      , (regs_regs_3_lpi_2[135:134]) , (regs_regs_3_lpi_2[137:136]) , (regs_regs_3_lpi_2[139:138])
      , (regs_regs_3_lpi_2[141:140]) , (regs_regs_3_lpi_2[143:142]) , (regs_regs_3_lpi_2[145:144])
      , (regs_regs_3_lpi_2[147:146]) , (regs_regs_3_lpi_2[149:148]) , (regs_regs_4_lpi_2[1:0])
      , (regs_regs_4_lpi_2[3:2]) , (regs_regs_4_lpi_2[5:4]) , (regs_regs_4_lpi_2[7:6])
      , (regs_regs_4_lpi_2[9:8]) , (regs_regs_4_lpi_2[11:10]) , (regs_regs_4_lpi_2[13:12])
      , (regs_regs_4_lpi_2[15:14]) , (regs_regs_4_lpi_2[17:16]) , (regs_regs_4_lpi_2[19:18])
      , (regs_regs_4_lpi_2[21:20]) , (regs_regs_4_lpi_2[23:22]) , (regs_regs_4_lpi_2[25:24])
      , (regs_regs_4_lpi_2[27:26]) , (regs_regs_4_lpi_2[29:28]) , (regs_regs_4_lpi_2[31:30])
      , (regs_regs_4_lpi_2[33:32]) , (regs_regs_4_lpi_2[35:34]) , (regs_regs_4_lpi_2[37:36])
      , (regs_regs_4_lpi_2[39:38]) , (regs_regs_4_lpi_2[41:40]) , (regs_regs_4_lpi_2[43:42])
      , (regs_regs_4_lpi_2[45:44]) , (regs_regs_4_lpi_2[47:46]) , (regs_regs_4_lpi_2[49:48])
      , (regs_regs_4_lpi_2[51:50]) , (regs_regs_4_lpi_2[53:52]) , (regs_regs_4_lpi_2[55:54])
      , (regs_regs_4_lpi_2[57:56]) , (regs_regs_4_lpi_2[59:58]) , (regs_regs_4_lpi_2[61:60])
      , (regs_regs_4_lpi_2[63:62]) , (regs_regs_4_lpi_2[65:64]) , (regs_regs_4_lpi_2[67:66])
      , (regs_regs_4_lpi_2[69:68]) , (regs_regs_4_lpi_2[71:70]) , (regs_regs_4_lpi_2[73:72])
      , (regs_regs_4_lpi_2[75:74]) , (regs_regs_4_lpi_2[77:76]) , (regs_regs_4_lpi_2[79:78])
      , (regs_regs_4_lpi_2[81:80]) , (regs_regs_4_lpi_2[83:82]) , (regs_regs_4_lpi_2[85:84])
      , (regs_regs_4_lpi_2[87:86]) , (regs_regs_4_lpi_2[89:88]) , (regs_regs_4_lpi_2[91:90])
      , (regs_regs_4_lpi_2[93:92]) , (regs_regs_4_lpi_2[95:94]) , (regs_regs_4_lpi_2[97:96])
      , (regs_regs_4_lpi_2[99:98]) , (regs_regs_4_lpi_2[101:100]) , (regs_regs_4_lpi_2[103:102])
      , (regs_regs_4_lpi_2[105:104]) , (regs_regs_4_lpi_2[107:106]) , (regs_regs_4_lpi_2[109:108])
      , (regs_regs_4_lpi_2[111:110]) , (regs_regs_4_lpi_2[113:112]) , (regs_regs_4_lpi_2[115:114])
      , (regs_regs_4_lpi_2[117:116]) , (regs_regs_4_lpi_2[119:118]) , (regs_regs_4_lpi_2[121:120])
      , (regs_regs_4_lpi_2[123:122]) , (regs_regs_4_lpi_2[125:124]) , (regs_regs_4_lpi_2[127:126])
      , (regs_regs_4_lpi_2[129:128]) , (regs_regs_4_lpi_2[131:130]) , (regs_regs_4_lpi_2[133:132])
      , (regs_regs_4_lpi_2[135:134]) , (regs_regs_4_lpi_2[137:136]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg7 = MUX_v_2_512_2({(regs_regs_0_lpi_2[15:14]) , (regs_regs_0_lpi_2[17:16])
      , (regs_regs_0_lpi_2[19:18]) , (regs_regs_0_lpi_2[21:20]) , (regs_regs_0_lpi_2[23:22])
      , (regs_regs_0_lpi_2[25:24]) , (regs_regs_0_lpi_2[27:26]) , (regs_regs_0_lpi_2[29:28])
      , (regs_regs_0_lpi_2[31:30]) , (regs_regs_0_lpi_2[33:32]) , (regs_regs_0_lpi_2[35:34])
      , (regs_regs_0_lpi_2[37:36]) , (regs_regs_0_lpi_2[39:38]) , (regs_regs_0_lpi_2[41:40])
      , (regs_regs_0_lpi_2[43:42]) , (regs_regs_0_lpi_2[45:44]) , (regs_regs_0_lpi_2[47:46])
      , (regs_regs_0_lpi_2[49:48]) , (regs_regs_0_lpi_2[51:50]) , (regs_regs_0_lpi_2[53:52])
      , (regs_regs_0_lpi_2[55:54]) , (regs_regs_0_lpi_2[57:56]) , (regs_regs_0_lpi_2[59:58])
      , (regs_regs_0_lpi_2[61:60]) , (regs_regs_0_lpi_2[63:62]) , (regs_regs_0_lpi_2[65:64])
      , (regs_regs_0_lpi_2[67:66]) , (regs_regs_0_lpi_2[69:68]) , (regs_regs_0_lpi_2[71:70])
      , (regs_regs_0_lpi_2[73:72]) , (regs_regs_0_lpi_2[75:74]) , (regs_regs_0_lpi_2[77:76])
      , (regs_regs_0_lpi_2[79:78]) , (regs_regs_0_lpi_2[81:80]) , (regs_regs_0_lpi_2[83:82])
      , (regs_regs_0_lpi_2[85:84]) , (regs_regs_0_lpi_2[87:86]) , (regs_regs_0_lpi_2[89:88])
      , (regs_regs_0_lpi_2[91:90]) , (regs_regs_0_lpi_2[93:92]) , (regs_regs_0_lpi_2[95:94])
      , (regs_regs_0_lpi_2[97:96]) , (regs_regs_0_lpi_2[99:98]) , (regs_regs_0_lpi_2[101:100])
      , (regs_regs_0_lpi_2[103:102]) , (regs_regs_0_lpi_2[105:104]) , (regs_regs_0_lpi_2[107:106])
      , (regs_regs_0_lpi_2[109:108]) , (regs_regs_0_lpi_2[111:110]) , (regs_regs_0_lpi_2[113:112])
      , (regs_regs_0_lpi_2[115:114]) , (regs_regs_0_lpi_2[117:116]) , (regs_regs_0_lpi_2[119:118])
      , (regs_regs_0_lpi_2[121:120]) , (regs_regs_0_lpi_2[123:122]) , (regs_regs_0_lpi_2[125:124])
      , (regs_regs_0_lpi_2[127:126]) , (regs_regs_0_lpi_2[129:128]) , (regs_regs_0_lpi_2[131:130])
      , (regs_regs_0_lpi_2[133:132]) , (regs_regs_0_lpi_2[135:134]) , (regs_regs_0_lpi_2[137:136])
      , (regs_regs_0_lpi_2[139:138]) , (regs_regs_0_lpi_2[141:140]) , (regs_regs_0_lpi_2[143:142])
      , (regs_regs_0_lpi_2[145:144]) , (regs_regs_0_lpi_2[147:146]) , (regs_regs_0_lpi_2[149:148])
      , (regs_regs_1_lpi_2[1:0]) , (regs_regs_1_lpi_2[3:2]) , (regs_regs_1_lpi_2[5:4])
      , (regs_regs_1_lpi_2[7:6]) , (regs_regs_1_lpi_2[9:8]) , (regs_regs_1_lpi_2[11:10])
      , (regs_regs_1_lpi_2[13:12]) , (regs_regs_1_lpi_2[15:14]) , (regs_regs_1_lpi_2[17:16])
      , (regs_regs_1_lpi_2[19:18]) , (regs_regs_1_lpi_2[21:20]) , (regs_regs_1_lpi_2[23:22])
      , (regs_regs_1_lpi_2[25:24]) , (regs_regs_1_lpi_2[27:26]) , (regs_regs_1_lpi_2[29:28])
      , (regs_regs_1_lpi_2[31:30]) , (regs_regs_1_lpi_2[33:32]) , (regs_regs_1_lpi_2[35:34])
      , (regs_regs_1_lpi_2[37:36]) , (regs_regs_1_lpi_2[39:38]) , (regs_regs_1_lpi_2[41:40])
      , (regs_regs_1_lpi_2[43:42]) , (regs_regs_1_lpi_2[45:44]) , (regs_regs_1_lpi_2[47:46])
      , (regs_regs_1_lpi_2[49:48]) , (regs_regs_1_lpi_2[51:50]) , (regs_regs_1_lpi_2[53:52])
      , (regs_regs_1_lpi_2[55:54]) , (regs_regs_1_lpi_2[57:56]) , (regs_regs_1_lpi_2[59:58])
      , (regs_regs_1_lpi_2[61:60]) , (regs_regs_1_lpi_2[63:62]) , (regs_regs_1_lpi_2[65:64])
      , (regs_regs_1_lpi_2[67:66]) , (regs_regs_1_lpi_2[69:68]) , (regs_regs_1_lpi_2[71:70])
      , (regs_regs_1_lpi_2[73:72]) , (regs_regs_1_lpi_2[75:74]) , (regs_regs_1_lpi_2[77:76])
      , (regs_regs_1_lpi_2[79:78]) , (regs_regs_1_lpi_2[81:80]) , (regs_regs_1_lpi_2[83:82])
      , (regs_regs_1_lpi_2[85:84]) , (regs_regs_1_lpi_2[87:86]) , (regs_regs_1_lpi_2[89:88])
      , (regs_regs_1_lpi_2[91:90]) , (regs_regs_1_lpi_2[93:92]) , (regs_regs_1_lpi_2[95:94])
      , (regs_regs_1_lpi_2[97:96]) , (regs_regs_1_lpi_2[99:98]) , (regs_regs_1_lpi_2[101:100])
      , (regs_regs_1_lpi_2[103:102]) , (regs_regs_1_lpi_2[105:104]) , (regs_regs_1_lpi_2[107:106])
      , (regs_regs_1_lpi_2[109:108]) , (regs_regs_1_lpi_2[111:110]) , (regs_regs_1_lpi_2[113:112])
      , (regs_regs_1_lpi_2[115:114]) , (regs_regs_1_lpi_2[117:116]) , (regs_regs_1_lpi_2[119:118])
      , (regs_regs_1_lpi_2[121:120]) , (regs_regs_1_lpi_2[123:122]) , (regs_regs_1_lpi_2[125:124])
      , (regs_regs_1_lpi_2[127:126]) , (regs_regs_1_lpi_2[129:128]) , (regs_regs_1_lpi_2[131:130])
      , (regs_regs_1_lpi_2[133:132]) , (regs_regs_1_lpi_2[135:134]) , (regs_regs_1_lpi_2[137:136])
      , (regs_regs_1_lpi_2[139:138]) , (regs_regs_1_lpi_2[141:140]) , (regs_regs_1_lpi_2[143:142])
      , (regs_regs_1_lpi_2[145:144]) , (regs_regs_1_lpi_2[147:146]) , (regs_regs_1_lpi_2[149:148])
      , (regs_regs_2_lpi_2[1:0]) , (regs_regs_2_lpi_2[3:2]) , (regs_regs_2_lpi_2[5:4])
      , (regs_regs_2_lpi_2[7:6]) , (regs_regs_2_lpi_2[9:8]) , (regs_regs_2_lpi_2[11:10])
      , (regs_regs_2_lpi_2[13:12]) , (regs_regs_2_lpi_2[15:14]) , (regs_regs_2_lpi_2[17:16])
      , (regs_regs_2_lpi_2[19:18]) , (regs_regs_2_lpi_2[21:20]) , (regs_regs_2_lpi_2[23:22])
      , (regs_regs_2_lpi_2[25:24]) , (regs_regs_2_lpi_2[27:26]) , (regs_regs_2_lpi_2[29:28])
      , (regs_regs_2_lpi_2[31:30]) , (regs_regs_2_lpi_2[33:32]) , (regs_regs_2_lpi_2[35:34])
      , (regs_regs_2_lpi_2[37:36]) , (regs_regs_2_lpi_2[39:38]) , (regs_regs_2_lpi_2[41:40])
      , (regs_regs_2_lpi_2[43:42]) , (regs_regs_2_lpi_2[45:44]) , (regs_regs_2_lpi_2[47:46])
      , (regs_regs_2_lpi_2[49:48]) , (regs_regs_2_lpi_2[51:50]) , (regs_regs_2_lpi_2[53:52])
      , (regs_regs_2_lpi_2[55:54]) , (regs_regs_2_lpi_2[57:56]) , (regs_regs_2_lpi_2[59:58])
      , (regs_regs_2_lpi_2[61:60]) , (regs_regs_2_lpi_2[63:62]) , (regs_regs_2_lpi_2[65:64])
      , (regs_regs_2_lpi_2[67:66]) , (regs_regs_2_lpi_2[69:68]) , (regs_regs_2_lpi_2[71:70])
      , (regs_regs_2_lpi_2[73:72]) , (regs_regs_2_lpi_2[75:74]) , (regs_regs_2_lpi_2[77:76])
      , (regs_regs_2_lpi_2[79:78]) , (regs_regs_2_lpi_2[81:80]) , (regs_regs_2_lpi_2[83:82])
      , (regs_regs_2_lpi_2[85:84]) , (regs_regs_2_lpi_2[87:86]) , (regs_regs_2_lpi_2[89:88])
      , (regs_regs_2_lpi_2[91:90]) , (regs_regs_2_lpi_2[93:92]) , (regs_regs_2_lpi_2[95:94])
      , (regs_regs_2_lpi_2[97:96]) , (regs_regs_2_lpi_2[99:98]) , (regs_regs_2_lpi_2[101:100])
      , (regs_regs_2_lpi_2[103:102]) , (regs_regs_2_lpi_2[105:104]) , (regs_regs_2_lpi_2[107:106])
      , (regs_regs_2_lpi_2[109:108]) , (regs_regs_2_lpi_2[111:110]) , (regs_regs_2_lpi_2[113:112])
      , (regs_regs_2_lpi_2[115:114]) , (regs_regs_2_lpi_2[117:116]) , (regs_regs_2_lpi_2[119:118])
      , (regs_regs_2_lpi_2[121:120]) , (regs_regs_2_lpi_2[123:122]) , (regs_regs_2_lpi_2[125:124])
      , (regs_regs_2_lpi_2[127:126]) , (regs_regs_2_lpi_2[129:128]) , (regs_regs_2_lpi_2[131:130])
      , (regs_regs_2_lpi_2[133:132]) , (regs_regs_2_lpi_2[135:134]) , (regs_regs_2_lpi_2[137:136])
      , (regs_regs_2_lpi_2[139:138]) , (regs_regs_2_lpi_2[141:140]) , (regs_regs_2_lpi_2[143:142])
      , (regs_regs_2_lpi_2[145:144]) , (regs_regs_2_lpi_2[147:146]) , (regs_regs_2_lpi_2[149:148])
      , (regs_regs_3_lpi_2[1:0]) , (regs_regs_3_lpi_2[3:2]) , (regs_regs_3_lpi_2[5:4])
      , (regs_regs_3_lpi_2[7:6]) , (regs_regs_3_lpi_2[9:8]) , (regs_regs_3_lpi_2[11:10])
      , (regs_regs_3_lpi_2[13:12]) , (regs_regs_3_lpi_2[15:14]) , (regs_regs_3_lpi_2[17:16])
      , (regs_regs_3_lpi_2[19:18]) , (regs_regs_3_lpi_2[21:20]) , (regs_regs_3_lpi_2[23:22])
      , (regs_regs_3_lpi_2[25:24]) , (regs_regs_3_lpi_2[27:26]) , (regs_regs_3_lpi_2[29:28])
      , (regs_regs_3_lpi_2[31:30]) , (regs_regs_3_lpi_2[33:32]) , (regs_regs_3_lpi_2[35:34])
      , (regs_regs_3_lpi_2[37:36]) , (regs_regs_3_lpi_2[39:38]) , (regs_regs_3_lpi_2[41:40])
      , (regs_regs_3_lpi_2[43:42]) , (regs_regs_3_lpi_2[45:44]) , (regs_regs_3_lpi_2[47:46])
      , (regs_regs_3_lpi_2[49:48]) , (regs_regs_3_lpi_2[51:50]) , (regs_regs_3_lpi_2[53:52])
      , (regs_regs_3_lpi_2[55:54]) , (regs_regs_3_lpi_2[57:56]) , (regs_regs_3_lpi_2[59:58])
      , (regs_regs_3_lpi_2[61:60]) , (regs_regs_3_lpi_2[63:62]) , (regs_regs_3_lpi_2[65:64])
      , (regs_regs_3_lpi_2[67:66]) , (regs_regs_3_lpi_2[69:68]) , (regs_regs_3_lpi_2[71:70])
      , (regs_regs_3_lpi_2[73:72]) , (regs_regs_3_lpi_2[75:74]) , (regs_regs_3_lpi_2[77:76])
      , (regs_regs_3_lpi_2[79:78]) , (regs_regs_3_lpi_2[81:80]) , (regs_regs_3_lpi_2[83:82])
      , (regs_regs_3_lpi_2[85:84]) , (regs_regs_3_lpi_2[87:86]) , (regs_regs_3_lpi_2[89:88])
      , (regs_regs_3_lpi_2[91:90]) , (regs_regs_3_lpi_2[93:92]) , (regs_regs_3_lpi_2[95:94])
      , (regs_regs_3_lpi_2[97:96]) , (regs_regs_3_lpi_2[99:98]) , (regs_regs_3_lpi_2[101:100])
      , (regs_regs_3_lpi_2[103:102]) , (regs_regs_3_lpi_2[105:104]) , (regs_regs_3_lpi_2[107:106])
      , (regs_regs_3_lpi_2[109:108]) , (regs_regs_3_lpi_2[111:110]) , (regs_regs_3_lpi_2[113:112])
      , (regs_regs_3_lpi_2[115:114]) , (regs_regs_3_lpi_2[117:116]) , (regs_regs_3_lpi_2[119:118])
      , (regs_regs_3_lpi_2[121:120]) , (regs_regs_3_lpi_2[123:122]) , (regs_regs_3_lpi_2[125:124])
      , (regs_regs_3_lpi_2[127:126]) , (regs_regs_3_lpi_2[129:128]) , (regs_regs_3_lpi_2[131:130])
      , (regs_regs_3_lpi_2[133:132]) , (regs_regs_3_lpi_2[135:134]) , (regs_regs_3_lpi_2[137:136])
      , (regs_regs_3_lpi_2[139:138]) , (regs_regs_3_lpi_2[141:140]) , (regs_regs_3_lpi_2[143:142])
      , (regs_regs_3_lpi_2[145:144]) , (regs_regs_3_lpi_2[147:146]) , (regs_regs_3_lpi_2[149:148])
      , (regs_regs_4_lpi_2[1:0]) , (regs_regs_4_lpi_2[3:2]) , (regs_regs_4_lpi_2[5:4])
      , (regs_regs_4_lpi_2[7:6]) , (regs_regs_4_lpi_2[9:8]) , (regs_regs_4_lpi_2[11:10])
      , (regs_regs_4_lpi_2[13:12]) , (regs_regs_4_lpi_2[15:14]) , (regs_regs_4_lpi_2[17:16])
      , (regs_regs_4_lpi_2[19:18]) , (regs_regs_4_lpi_2[21:20]) , (regs_regs_4_lpi_2[23:22])
      , (regs_regs_4_lpi_2[25:24]) , (regs_regs_4_lpi_2[27:26]) , (regs_regs_4_lpi_2[29:28])
      , (regs_regs_4_lpi_2[31:30]) , (regs_regs_4_lpi_2[33:32]) , (regs_regs_4_lpi_2[35:34])
      , (regs_regs_4_lpi_2[37:36]) , (regs_regs_4_lpi_2[39:38]) , (regs_regs_4_lpi_2[41:40])
      , (regs_regs_4_lpi_2[43:42]) , (regs_regs_4_lpi_2[45:44]) , (regs_regs_4_lpi_2[47:46])
      , (regs_regs_4_lpi_2[49:48]) , (regs_regs_4_lpi_2[51:50]) , (regs_regs_4_lpi_2[53:52])
      , (regs_regs_4_lpi_2[55:54]) , (regs_regs_4_lpi_2[57:56]) , (regs_regs_4_lpi_2[59:58])
      , (regs_regs_4_lpi_2[61:60]) , (regs_regs_4_lpi_2[63:62]) , (regs_regs_4_lpi_2[65:64])
      , (regs_regs_4_lpi_2[67:66]) , (regs_regs_4_lpi_2[69:68]) , (regs_regs_4_lpi_2[71:70])
      , (regs_regs_4_lpi_2[73:72]) , (regs_regs_4_lpi_2[75:74]) , (regs_regs_4_lpi_2[77:76])
      , (regs_regs_4_lpi_2[79:78]) , (regs_regs_4_lpi_2[81:80]) , (regs_regs_4_lpi_2[83:82])
      , (regs_regs_4_lpi_2[85:84]) , (regs_regs_4_lpi_2[87:86]) , (regs_regs_4_lpi_2[89:88])
      , (regs_regs_4_lpi_2[91:90]) , (regs_regs_4_lpi_2[93:92]) , (regs_regs_4_lpi_2[95:94])
      , (regs_regs_4_lpi_2[97:96]) , (regs_regs_4_lpi_2[99:98]) , (regs_regs_4_lpi_2[101:100])
      , (regs_regs_4_lpi_2[103:102]) , (regs_regs_4_lpi_2[105:104]) , (regs_regs_4_lpi_2[107:106])
      , (regs_regs_4_lpi_2[109:108]) , (regs_regs_4_lpi_2[111:110]) , (regs_regs_4_lpi_2[113:112])
      , (regs_regs_4_lpi_2[115:114]) , (regs_regs_4_lpi_2[117:116]) , (regs_regs_4_lpi_2[119:118])
      , (regs_regs_4_lpi_2[121:120]) , (regs_regs_4_lpi_2[123:122]) , (regs_regs_4_lpi_2[125:124])
      , (regs_regs_4_lpi_2[127:126]) , (regs_regs_4_lpi_2[129:128]) , (regs_regs_4_lpi_2[131:130])
      , (regs_regs_4_lpi_2[133:132]) , (regs_regs_4_lpi_2[135:134]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg6 = MUX_v_2_512_2({(regs_regs_0_lpi_2[13:12]) , (regs_regs_0_lpi_2[15:14])
      , (regs_regs_0_lpi_2[17:16]) , (regs_regs_0_lpi_2[19:18]) , (regs_regs_0_lpi_2[21:20])
      , (regs_regs_0_lpi_2[23:22]) , (regs_regs_0_lpi_2[25:24]) , (regs_regs_0_lpi_2[27:26])
      , (regs_regs_0_lpi_2[29:28]) , (regs_regs_0_lpi_2[31:30]) , (regs_regs_0_lpi_2[33:32])
      , (regs_regs_0_lpi_2[35:34]) , (regs_regs_0_lpi_2[37:36]) , (regs_regs_0_lpi_2[39:38])
      , (regs_regs_0_lpi_2[41:40]) , (regs_regs_0_lpi_2[43:42]) , (regs_regs_0_lpi_2[45:44])
      , (regs_regs_0_lpi_2[47:46]) , (regs_regs_0_lpi_2[49:48]) , (regs_regs_0_lpi_2[51:50])
      , (regs_regs_0_lpi_2[53:52]) , (regs_regs_0_lpi_2[55:54]) , (regs_regs_0_lpi_2[57:56])
      , (regs_regs_0_lpi_2[59:58]) , (regs_regs_0_lpi_2[61:60]) , (regs_regs_0_lpi_2[63:62])
      , (regs_regs_0_lpi_2[65:64]) , (regs_regs_0_lpi_2[67:66]) , (regs_regs_0_lpi_2[69:68])
      , (regs_regs_0_lpi_2[71:70]) , (regs_regs_0_lpi_2[73:72]) , (regs_regs_0_lpi_2[75:74])
      , (regs_regs_0_lpi_2[77:76]) , (regs_regs_0_lpi_2[79:78]) , (regs_regs_0_lpi_2[81:80])
      , (regs_regs_0_lpi_2[83:82]) , (regs_regs_0_lpi_2[85:84]) , (regs_regs_0_lpi_2[87:86])
      , (regs_regs_0_lpi_2[89:88]) , (regs_regs_0_lpi_2[91:90]) , (regs_regs_0_lpi_2[93:92])
      , (regs_regs_0_lpi_2[95:94]) , (regs_regs_0_lpi_2[97:96]) , (regs_regs_0_lpi_2[99:98])
      , (regs_regs_0_lpi_2[101:100]) , (regs_regs_0_lpi_2[103:102]) , (regs_regs_0_lpi_2[105:104])
      , (regs_regs_0_lpi_2[107:106]) , (regs_regs_0_lpi_2[109:108]) , (regs_regs_0_lpi_2[111:110])
      , (regs_regs_0_lpi_2[113:112]) , (regs_regs_0_lpi_2[115:114]) , (regs_regs_0_lpi_2[117:116])
      , (regs_regs_0_lpi_2[119:118]) , (regs_regs_0_lpi_2[121:120]) , (regs_regs_0_lpi_2[123:122])
      , (regs_regs_0_lpi_2[125:124]) , (regs_regs_0_lpi_2[127:126]) , (regs_regs_0_lpi_2[129:128])
      , (regs_regs_0_lpi_2[131:130]) , (regs_regs_0_lpi_2[133:132]) , (regs_regs_0_lpi_2[135:134])
      , (regs_regs_0_lpi_2[137:136]) , (regs_regs_0_lpi_2[139:138]) , (regs_regs_0_lpi_2[141:140])
      , (regs_regs_0_lpi_2[143:142]) , (regs_regs_0_lpi_2[145:144]) , (regs_regs_0_lpi_2[147:146])
      , (regs_regs_0_lpi_2[149:148]) , (regs_regs_1_lpi_2[1:0]) , (regs_regs_1_lpi_2[3:2])
      , (regs_regs_1_lpi_2[5:4]) , (regs_regs_1_lpi_2[7:6]) , (regs_regs_1_lpi_2[9:8])
      , (regs_regs_1_lpi_2[11:10]) , (regs_regs_1_lpi_2[13:12]) , (regs_regs_1_lpi_2[15:14])
      , (regs_regs_1_lpi_2[17:16]) , (regs_regs_1_lpi_2[19:18]) , (regs_regs_1_lpi_2[21:20])
      , (regs_regs_1_lpi_2[23:22]) , (regs_regs_1_lpi_2[25:24]) , (regs_regs_1_lpi_2[27:26])
      , (regs_regs_1_lpi_2[29:28]) , (regs_regs_1_lpi_2[31:30]) , (regs_regs_1_lpi_2[33:32])
      , (regs_regs_1_lpi_2[35:34]) , (regs_regs_1_lpi_2[37:36]) , (regs_regs_1_lpi_2[39:38])
      , (regs_regs_1_lpi_2[41:40]) , (regs_regs_1_lpi_2[43:42]) , (regs_regs_1_lpi_2[45:44])
      , (regs_regs_1_lpi_2[47:46]) , (regs_regs_1_lpi_2[49:48]) , (regs_regs_1_lpi_2[51:50])
      , (regs_regs_1_lpi_2[53:52]) , (regs_regs_1_lpi_2[55:54]) , (regs_regs_1_lpi_2[57:56])
      , (regs_regs_1_lpi_2[59:58]) , (regs_regs_1_lpi_2[61:60]) , (regs_regs_1_lpi_2[63:62])
      , (regs_regs_1_lpi_2[65:64]) , (regs_regs_1_lpi_2[67:66]) , (regs_regs_1_lpi_2[69:68])
      , (regs_regs_1_lpi_2[71:70]) , (regs_regs_1_lpi_2[73:72]) , (regs_regs_1_lpi_2[75:74])
      , (regs_regs_1_lpi_2[77:76]) , (regs_regs_1_lpi_2[79:78]) , (regs_regs_1_lpi_2[81:80])
      , (regs_regs_1_lpi_2[83:82]) , (regs_regs_1_lpi_2[85:84]) , (regs_regs_1_lpi_2[87:86])
      , (regs_regs_1_lpi_2[89:88]) , (regs_regs_1_lpi_2[91:90]) , (regs_regs_1_lpi_2[93:92])
      , (regs_regs_1_lpi_2[95:94]) , (regs_regs_1_lpi_2[97:96]) , (regs_regs_1_lpi_2[99:98])
      , (regs_regs_1_lpi_2[101:100]) , (regs_regs_1_lpi_2[103:102]) , (regs_regs_1_lpi_2[105:104])
      , (regs_regs_1_lpi_2[107:106]) , (regs_regs_1_lpi_2[109:108]) , (regs_regs_1_lpi_2[111:110])
      , (regs_regs_1_lpi_2[113:112]) , (regs_regs_1_lpi_2[115:114]) , (regs_regs_1_lpi_2[117:116])
      , (regs_regs_1_lpi_2[119:118]) , (regs_regs_1_lpi_2[121:120]) , (regs_regs_1_lpi_2[123:122])
      , (regs_regs_1_lpi_2[125:124]) , (regs_regs_1_lpi_2[127:126]) , (regs_regs_1_lpi_2[129:128])
      , (regs_regs_1_lpi_2[131:130]) , (regs_regs_1_lpi_2[133:132]) , (regs_regs_1_lpi_2[135:134])
      , (regs_regs_1_lpi_2[137:136]) , (regs_regs_1_lpi_2[139:138]) , (regs_regs_1_lpi_2[141:140])
      , (regs_regs_1_lpi_2[143:142]) , (regs_regs_1_lpi_2[145:144]) , (regs_regs_1_lpi_2[147:146])
      , (regs_regs_1_lpi_2[149:148]) , (regs_regs_2_lpi_2[1:0]) , (regs_regs_2_lpi_2[3:2])
      , (regs_regs_2_lpi_2[5:4]) , (regs_regs_2_lpi_2[7:6]) , (regs_regs_2_lpi_2[9:8])
      , (regs_regs_2_lpi_2[11:10]) , (regs_regs_2_lpi_2[13:12]) , (regs_regs_2_lpi_2[15:14])
      , (regs_regs_2_lpi_2[17:16]) , (regs_regs_2_lpi_2[19:18]) , (regs_regs_2_lpi_2[21:20])
      , (regs_regs_2_lpi_2[23:22]) , (regs_regs_2_lpi_2[25:24]) , (regs_regs_2_lpi_2[27:26])
      , (regs_regs_2_lpi_2[29:28]) , (regs_regs_2_lpi_2[31:30]) , (regs_regs_2_lpi_2[33:32])
      , (regs_regs_2_lpi_2[35:34]) , (regs_regs_2_lpi_2[37:36]) , (regs_regs_2_lpi_2[39:38])
      , (regs_regs_2_lpi_2[41:40]) , (regs_regs_2_lpi_2[43:42]) , (regs_regs_2_lpi_2[45:44])
      , (regs_regs_2_lpi_2[47:46]) , (regs_regs_2_lpi_2[49:48]) , (regs_regs_2_lpi_2[51:50])
      , (regs_regs_2_lpi_2[53:52]) , (regs_regs_2_lpi_2[55:54]) , (regs_regs_2_lpi_2[57:56])
      , (regs_regs_2_lpi_2[59:58]) , (regs_regs_2_lpi_2[61:60]) , (regs_regs_2_lpi_2[63:62])
      , (regs_regs_2_lpi_2[65:64]) , (regs_regs_2_lpi_2[67:66]) , (regs_regs_2_lpi_2[69:68])
      , (regs_regs_2_lpi_2[71:70]) , (regs_regs_2_lpi_2[73:72]) , (regs_regs_2_lpi_2[75:74])
      , (regs_regs_2_lpi_2[77:76]) , (regs_regs_2_lpi_2[79:78]) , (regs_regs_2_lpi_2[81:80])
      , (regs_regs_2_lpi_2[83:82]) , (regs_regs_2_lpi_2[85:84]) , (regs_regs_2_lpi_2[87:86])
      , (regs_regs_2_lpi_2[89:88]) , (regs_regs_2_lpi_2[91:90]) , (regs_regs_2_lpi_2[93:92])
      , (regs_regs_2_lpi_2[95:94]) , (regs_regs_2_lpi_2[97:96]) , (regs_regs_2_lpi_2[99:98])
      , (regs_regs_2_lpi_2[101:100]) , (regs_regs_2_lpi_2[103:102]) , (regs_regs_2_lpi_2[105:104])
      , (regs_regs_2_lpi_2[107:106]) , (regs_regs_2_lpi_2[109:108]) , (regs_regs_2_lpi_2[111:110])
      , (regs_regs_2_lpi_2[113:112]) , (regs_regs_2_lpi_2[115:114]) , (regs_regs_2_lpi_2[117:116])
      , (regs_regs_2_lpi_2[119:118]) , (regs_regs_2_lpi_2[121:120]) , (regs_regs_2_lpi_2[123:122])
      , (regs_regs_2_lpi_2[125:124]) , (regs_regs_2_lpi_2[127:126]) , (regs_regs_2_lpi_2[129:128])
      , (regs_regs_2_lpi_2[131:130]) , (regs_regs_2_lpi_2[133:132]) , (regs_regs_2_lpi_2[135:134])
      , (regs_regs_2_lpi_2[137:136]) , (regs_regs_2_lpi_2[139:138]) , (regs_regs_2_lpi_2[141:140])
      , (regs_regs_2_lpi_2[143:142]) , (regs_regs_2_lpi_2[145:144]) , (regs_regs_2_lpi_2[147:146])
      , (regs_regs_2_lpi_2[149:148]) , (regs_regs_3_lpi_2[1:0]) , (regs_regs_3_lpi_2[3:2])
      , (regs_regs_3_lpi_2[5:4]) , (regs_regs_3_lpi_2[7:6]) , (regs_regs_3_lpi_2[9:8])
      , (regs_regs_3_lpi_2[11:10]) , (regs_regs_3_lpi_2[13:12]) , (regs_regs_3_lpi_2[15:14])
      , (regs_regs_3_lpi_2[17:16]) , (regs_regs_3_lpi_2[19:18]) , (regs_regs_3_lpi_2[21:20])
      , (regs_regs_3_lpi_2[23:22]) , (regs_regs_3_lpi_2[25:24]) , (regs_regs_3_lpi_2[27:26])
      , (regs_regs_3_lpi_2[29:28]) , (regs_regs_3_lpi_2[31:30]) , (regs_regs_3_lpi_2[33:32])
      , (regs_regs_3_lpi_2[35:34]) , (regs_regs_3_lpi_2[37:36]) , (regs_regs_3_lpi_2[39:38])
      , (regs_regs_3_lpi_2[41:40]) , (regs_regs_3_lpi_2[43:42]) , (regs_regs_3_lpi_2[45:44])
      , (regs_regs_3_lpi_2[47:46]) , (regs_regs_3_lpi_2[49:48]) , (regs_regs_3_lpi_2[51:50])
      , (regs_regs_3_lpi_2[53:52]) , (regs_regs_3_lpi_2[55:54]) , (regs_regs_3_lpi_2[57:56])
      , (regs_regs_3_lpi_2[59:58]) , (regs_regs_3_lpi_2[61:60]) , (regs_regs_3_lpi_2[63:62])
      , (regs_regs_3_lpi_2[65:64]) , (regs_regs_3_lpi_2[67:66]) , (regs_regs_3_lpi_2[69:68])
      , (regs_regs_3_lpi_2[71:70]) , (regs_regs_3_lpi_2[73:72]) , (regs_regs_3_lpi_2[75:74])
      , (regs_regs_3_lpi_2[77:76]) , (regs_regs_3_lpi_2[79:78]) , (regs_regs_3_lpi_2[81:80])
      , (regs_regs_3_lpi_2[83:82]) , (regs_regs_3_lpi_2[85:84]) , (regs_regs_3_lpi_2[87:86])
      , (regs_regs_3_lpi_2[89:88]) , (regs_regs_3_lpi_2[91:90]) , (regs_regs_3_lpi_2[93:92])
      , (regs_regs_3_lpi_2[95:94]) , (regs_regs_3_lpi_2[97:96]) , (regs_regs_3_lpi_2[99:98])
      , (regs_regs_3_lpi_2[101:100]) , (regs_regs_3_lpi_2[103:102]) , (regs_regs_3_lpi_2[105:104])
      , (regs_regs_3_lpi_2[107:106]) , (regs_regs_3_lpi_2[109:108]) , (regs_regs_3_lpi_2[111:110])
      , (regs_regs_3_lpi_2[113:112]) , (regs_regs_3_lpi_2[115:114]) , (regs_regs_3_lpi_2[117:116])
      , (regs_regs_3_lpi_2[119:118]) , (regs_regs_3_lpi_2[121:120]) , (regs_regs_3_lpi_2[123:122])
      , (regs_regs_3_lpi_2[125:124]) , (regs_regs_3_lpi_2[127:126]) , (regs_regs_3_lpi_2[129:128])
      , (regs_regs_3_lpi_2[131:130]) , (regs_regs_3_lpi_2[133:132]) , (regs_regs_3_lpi_2[135:134])
      , (regs_regs_3_lpi_2[137:136]) , (regs_regs_3_lpi_2[139:138]) , (regs_regs_3_lpi_2[141:140])
      , (regs_regs_3_lpi_2[143:142]) , (regs_regs_3_lpi_2[145:144]) , (regs_regs_3_lpi_2[147:146])
      , (regs_regs_3_lpi_2[149:148]) , (regs_regs_4_lpi_2[1:0]) , (regs_regs_4_lpi_2[3:2])
      , (regs_regs_4_lpi_2[5:4]) , (regs_regs_4_lpi_2[7:6]) , (regs_regs_4_lpi_2[9:8])
      , (regs_regs_4_lpi_2[11:10]) , (regs_regs_4_lpi_2[13:12]) , (regs_regs_4_lpi_2[15:14])
      , (regs_regs_4_lpi_2[17:16]) , (regs_regs_4_lpi_2[19:18]) , (regs_regs_4_lpi_2[21:20])
      , (regs_regs_4_lpi_2[23:22]) , (regs_regs_4_lpi_2[25:24]) , (regs_regs_4_lpi_2[27:26])
      , (regs_regs_4_lpi_2[29:28]) , (regs_regs_4_lpi_2[31:30]) , (regs_regs_4_lpi_2[33:32])
      , (regs_regs_4_lpi_2[35:34]) , (regs_regs_4_lpi_2[37:36]) , (regs_regs_4_lpi_2[39:38])
      , (regs_regs_4_lpi_2[41:40]) , (regs_regs_4_lpi_2[43:42]) , (regs_regs_4_lpi_2[45:44])
      , (regs_regs_4_lpi_2[47:46]) , (regs_regs_4_lpi_2[49:48]) , (regs_regs_4_lpi_2[51:50])
      , (regs_regs_4_lpi_2[53:52]) , (regs_regs_4_lpi_2[55:54]) , (regs_regs_4_lpi_2[57:56])
      , (regs_regs_4_lpi_2[59:58]) , (regs_regs_4_lpi_2[61:60]) , (regs_regs_4_lpi_2[63:62])
      , (regs_regs_4_lpi_2[65:64]) , (regs_regs_4_lpi_2[67:66]) , (regs_regs_4_lpi_2[69:68])
      , (regs_regs_4_lpi_2[71:70]) , (regs_regs_4_lpi_2[73:72]) , (regs_regs_4_lpi_2[75:74])
      , (regs_regs_4_lpi_2[77:76]) , (regs_regs_4_lpi_2[79:78]) , (regs_regs_4_lpi_2[81:80])
      , (regs_regs_4_lpi_2[83:82]) , (regs_regs_4_lpi_2[85:84]) , (regs_regs_4_lpi_2[87:86])
      , (regs_regs_4_lpi_2[89:88]) , (regs_regs_4_lpi_2[91:90]) , (regs_regs_4_lpi_2[93:92])
      , (regs_regs_4_lpi_2[95:94]) , (regs_regs_4_lpi_2[97:96]) , (regs_regs_4_lpi_2[99:98])
      , (regs_regs_4_lpi_2[101:100]) , (regs_regs_4_lpi_2[103:102]) , (regs_regs_4_lpi_2[105:104])
      , (regs_regs_4_lpi_2[107:106]) , (regs_regs_4_lpi_2[109:108]) , (regs_regs_4_lpi_2[111:110])
      , (regs_regs_4_lpi_2[113:112]) , (regs_regs_4_lpi_2[115:114]) , (regs_regs_4_lpi_2[117:116])
      , (regs_regs_4_lpi_2[119:118]) , (regs_regs_4_lpi_2[121:120]) , (regs_regs_4_lpi_2[123:122])
      , (regs_regs_4_lpi_2[125:124]) , (regs_regs_4_lpi_2[127:126]) , (regs_regs_4_lpi_2[129:128])
      , (regs_regs_4_lpi_2[131:130]) , (regs_regs_4_lpi_2[133:132]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg5 = MUX_v_2_512_2({(regs_regs_0_lpi_2[11:10]) , (regs_regs_0_lpi_2[13:12])
      , (regs_regs_0_lpi_2[15:14]) , (regs_regs_0_lpi_2[17:16]) , (regs_regs_0_lpi_2[19:18])
      , (regs_regs_0_lpi_2[21:20]) , (regs_regs_0_lpi_2[23:22]) , (regs_regs_0_lpi_2[25:24])
      , (regs_regs_0_lpi_2[27:26]) , (regs_regs_0_lpi_2[29:28]) , (regs_regs_0_lpi_2[31:30])
      , (regs_regs_0_lpi_2[33:32]) , (regs_regs_0_lpi_2[35:34]) , (regs_regs_0_lpi_2[37:36])
      , (regs_regs_0_lpi_2[39:38]) , (regs_regs_0_lpi_2[41:40]) , (regs_regs_0_lpi_2[43:42])
      , (regs_regs_0_lpi_2[45:44]) , (regs_regs_0_lpi_2[47:46]) , (regs_regs_0_lpi_2[49:48])
      , (regs_regs_0_lpi_2[51:50]) , (regs_regs_0_lpi_2[53:52]) , (regs_regs_0_lpi_2[55:54])
      , (regs_regs_0_lpi_2[57:56]) , (regs_regs_0_lpi_2[59:58]) , (regs_regs_0_lpi_2[61:60])
      , (regs_regs_0_lpi_2[63:62]) , (regs_regs_0_lpi_2[65:64]) , (regs_regs_0_lpi_2[67:66])
      , (regs_regs_0_lpi_2[69:68]) , (regs_regs_0_lpi_2[71:70]) , (regs_regs_0_lpi_2[73:72])
      , (regs_regs_0_lpi_2[75:74]) , (regs_regs_0_lpi_2[77:76]) , (regs_regs_0_lpi_2[79:78])
      , (regs_regs_0_lpi_2[81:80]) , (regs_regs_0_lpi_2[83:82]) , (regs_regs_0_lpi_2[85:84])
      , (regs_regs_0_lpi_2[87:86]) , (regs_regs_0_lpi_2[89:88]) , (regs_regs_0_lpi_2[91:90])
      , (regs_regs_0_lpi_2[93:92]) , (regs_regs_0_lpi_2[95:94]) , (regs_regs_0_lpi_2[97:96])
      , (regs_regs_0_lpi_2[99:98]) , (regs_regs_0_lpi_2[101:100]) , (regs_regs_0_lpi_2[103:102])
      , (regs_regs_0_lpi_2[105:104]) , (regs_regs_0_lpi_2[107:106]) , (regs_regs_0_lpi_2[109:108])
      , (regs_regs_0_lpi_2[111:110]) , (regs_regs_0_lpi_2[113:112]) , (regs_regs_0_lpi_2[115:114])
      , (regs_regs_0_lpi_2[117:116]) , (regs_regs_0_lpi_2[119:118]) , (regs_regs_0_lpi_2[121:120])
      , (regs_regs_0_lpi_2[123:122]) , (regs_regs_0_lpi_2[125:124]) , (regs_regs_0_lpi_2[127:126])
      , (regs_regs_0_lpi_2[129:128]) , (regs_regs_0_lpi_2[131:130]) , (regs_regs_0_lpi_2[133:132])
      , (regs_regs_0_lpi_2[135:134]) , (regs_regs_0_lpi_2[137:136]) , (regs_regs_0_lpi_2[139:138])
      , (regs_regs_0_lpi_2[141:140]) , (regs_regs_0_lpi_2[143:142]) , (regs_regs_0_lpi_2[145:144])
      , (regs_regs_0_lpi_2[147:146]) , (regs_regs_0_lpi_2[149:148]) , (regs_regs_1_lpi_2[1:0])
      , (regs_regs_1_lpi_2[3:2]) , (regs_regs_1_lpi_2[5:4]) , (regs_regs_1_lpi_2[7:6])
      , (regs_regs_1_lpi_2[9:8]) , (regs_regs_1_lpi_2[11:10]) , (regs_regs_1_lpi_2[13:12])
      , (regs_regs_1_lpi_2[15:14]) , (regs_regs_1_lpi_2[17:16]) , (regs_regs_1_lpi_2[19:18])
      , (regs_regs_1_lpi_2[21:20]) , (regs_regs_1_lpi_2[23:22]) , (regs_regs_1_lpi_2[25:24])
      , (regs_regs_1_lpi_2[27:26]) , (regs_regs_1_lpi_2[29:28]) , (regs_regs_1_lpi_2[31:30])
      , (regs_regs_1_lpi_2[33:32]) , (regs_regs_1_lpi_2[35:34]) , (regs_regs_1_lpi_2[37:36])
      , (regs_regs_1_lpi_2[39:38]) , (regs_regs_1_lpi_2[41:40]) , (regs_regs_1_lpi_2[43:42])
      , (regs_regs_1_lpi_2[45:44]) , (regs_regs_1_lpi_2[47:46]) , (regs_regs_1_lpi_2[49:48])
      , (regs_regs_1_lpi_2[51:50]) , (regs_regs_1_lpi_2[53:52]) , (regs_regs_1_lpi_2[55:54])
      , (regs_regs_1_lpi_2[57:56]) , (regs_regs_1_lpi_2[59:58]) , (regs_regs_1_lpi_2[61:60])
      , (regs_regs_1_lpi_2[63:62]) , (regs_regs_1_lpi_2[65:64]) , (regs_regs_1_lpi_2[67:66])
      , (regs_regs_1_lpi_2[69:68]) , (regs_regs_1_lpi_2[71:70]) , (regs_regs_1_lpi_2[73:72])
      , (regs_regs_1_lpi_2[75:74]) , (regs_regs_1_lpi_2[77:76]) , (regs_regs_1_lpi_2[79:78])
      , (regs_regs_1_lpi_2[81:80]) , (regs_regs_1_lpi_2[83:82]) , (regs_regs_1_lpi_2[85:84])
      , (regs_regs_1_lpi_2[87:86]) , (regs_regs_1_lpi_2[89:88]) , (regs_regs_1_lpi_2[91:90])
      , (regs_regs_1_lpi_2[93:92]) , (regs_regs_1_lpi_2[95:94]) , (regs_regs_1_lpi_2[97:96])
      , (regs_regs_1_lpi_2[99:98]) , (regs_regs_1_lpi_2[101:100]) , (regs_regs_1_lpi_2[103:102])
      , (regs_regs_1_lpi_2[105:104]) , (regs_regs_1_lpi_2[107:106]) , (regs_regs_1_lpi_2[109:108])
      , (regs_regs_1_lpi_2[111:110]) , (regs_regs_1_lpi_2[113:112]) , (regs_regs_1_lpi_2[115:114])
      , (regs_regs_1_lpi_2[117:116]) , (regs_regs_1_lpi_2[119:118]) , (regs_regs_1_lpi_2[121:120])
      , (regs_regs_1_lpi_2[123:122]) , (regs_regs_1_lpi_2[125:124]) , (regs_regs_1_lpi_2[127:126])
      , (regs_regs_1_lpi_2[129:128]) , (regs_regs_1_lpi_2[131:130]) , (regs_regs_1_lpi_2[133:132])
      , (regs_regs_1_lpi_2[135:134]) , (regs_regs_1_lpi_2[137:136]) , (regs_regs_1_lpi_2[139:138])
      , (regs_regs_1_lpi_2[141:140]) , (regs_regs_1_lpi_2[143:142]) , (regs_regs_1_lpi_2[145:144])
      , (regs_regs_1_lpi_2[147:146]) , (regs_regs_1_lpi_2[149:148]) , (regs_regs_2_lpi_2[1:0])
      , (regs_regs_2_lpi_2[3:2]) , (regs_regs_2_lpi_2[5:4]) , (regs_regs_2_lpi_2[7:6])
      , (regs_regs_2_lpi_2[9:8]) , (regs_regs_2_lpi_2[11:10]) , (regs_regs_2_lpi_2[13:12])
      , (regs_regs_2_lpi_2[15:14]) , (regs_regs_2_lpi_2[17:16]) , (regs_regs_2_lpi_2[19:18])
      , (regs_regs_2_lpi_2[21:20]) , (regs_regs_2_lpi_2[23:22]) , (regs_regs_2_lpi_2[25:24])
      , (regs_regs_2_lpi_2[27:26]) , (regs_regs_2_lpi_2[29:28]) , (regs_regs_2_lpi_2[31:30])
      , (regs_regs_2_lpi_2[33:32]) , (regs_regs_2_lpi_2[35:34]) , (regs_regs_2_lpi_2[37:36])
      , (regs_regs_2_lpi_2[39:38]) , (regs_regs_2_lpi_2[41:40]) , (regs_regs_2_lpi_2[43:42])
      , (regs_regs_2_lpi_2[45:44]) , (regs_regs_2_lpi_2[47:46]) , (regs_regs_2_lpi_2[49:48])
      , (regs_regs_2_lpi_2[51:50]) , (regs_regs_2_lpi_2[53:52]) , (regs_regs_2_lpi_2[55:54])
      , (regs_regs_2_lpi_2[57:56]) , (regs_regs_2_lpi_2[59:58]) , (regs_regs_2_lpi_2[61:60])
      , (regs_regs_2_lpi_2[63:62]) , (regs_regs_2_lpi_2[65:64]) , (regs_regs_2_lpi_2[67:66])
      , (regs_regs_2_lpi_2[69:68]) , (regs_regs_2_lpi_2[71:70]) , (regs_regs_2_lpi_2[73:72])
      , (regs_regs_2_lpi_2[75:74]) , (regs_regs_2_lpi_2[77:76]) , (regs_regs_2_lpi_2[79:78])
      , (regs_regs_2_lpi_2[81:80]) , (regs_regs_2_lpi_2[83:82]) , (regs_regs_2_lpi_2[85:84])
      , (regs_regs_2_lpi_2[87:86]) , (regs_regs_2_lpi_2[89:88]) , (regs_regs_2_lpi_2[91:90])
      , (regs_regs_2_lpi_2[93:92]) , (regs_regs_2_lpi_2[95:94]) , (regs_regs_2_lpi_2[97:96])
      , (regs_regs_2_lpi_2[99:98]) , (regs_regs_2_lpi_2[101:100]) , (regs_regs_2_lpi_2[103:102])
      , (regs_regs_2_lpi_2[105:104]) , (regs_regs_2_lpi_2[107:106]) , (regs_regs_2_lpi_2[109:108])
      , (regs_regs_2_lpi_2[111:110]) , (regs_regs_2_lpi_2[113:112]) , (regs_regs_2_lpi_2[115:114])
      , (regs_regs_2_lpi_2[117:116]) , (regs_regs_2_lpi_2[119:118]) , (regs_regs_2_lpi_2[121:120])
      , (regs_regs_2_lpi_2[123:122]) , (regs_regs_2_lpi_2[125:124]) , (regs_regs_2_lpi_2[127:126])
      , (regs_regs_2_lpi_2[129:128]) , (regs_regs_2_lpi_2[131:130]) , (regs_regs_2_lpi_2[133:132])
      , (regs_regs_2_lpi_2[135:134]) , (regs_regs_2_lpi_2[137:136]) , (regs_regs_2_lpi_2[139:138])
      , (regs_regs_2_lpi_2[141:140]) , (regs_regs_2_lpi_2[143:142]) , (regs_regs_2_lpi_2[145:144])
      , (regs_regs_2_lpi_2[147:146]) , (regs_regs_2_lpi_2[149:148]) , (regs_regs_3_lpi_2[1:0])
      , (regs_regs_3_lpi_2[3:2]) , (regs_regs_3_lpi_2[5:4]) , (regs_regs_3_lpi_2[7:6])
      , (regs_regs_3_lpi_2[9:8]) , (regs_regs_3_lpi_2[11:10]) , (regs_regs_3_lpi_2[13:12])
      , (regs_regs_3_lpi_2[15:14]) , (regs_regs_3_lpi_2[17:16]) , (regs_regs_3_lpi_2[19:18])
      , (regs_regs_3_lpi_2[21:20]) , (regs_regs_3_lpi_2[23:22]) , (regs_regs_3_lpi_2[25:24])
      , (regs_regs_3_lpi_2[27:26]) , (regs_regs_3_lpi_2[29:28]) , (regs_regs_3_lpi_2[31:30])
      , (regs_regs_3_lpi_2[33:32]) , (regs_regs_3_lpi_2[35:34]) , (regs_regs_3_lpi_2[37:36])
      , (regs_regs_3_lpi_2[39:38]) , (regs_regs_3_lpi_2[41:40]) , (regs_regs_3_lpi_2[43:42])
      , (regs_regs_3_lpi_2[45:44]) , (regs_regs_3_lpi_2[47:46]) , (regs_regs_3_lpi_2[49:48])
      , (regs_regs_3_lpi_2[51:50]) , (regs_regs_3_lpi_2[53:52]) , (regs_regs_3_lpi_2[55:54])
      , (regs_regs_3_lpi_2[57:56]) , (regs_regs_3_lpi_2[59:58]) , (regs_regs_3_lpi_2[61:60])
      , (regs_regs_3_lpi_2[63:62]) , (regs_regs_3_lpi_2[65:64]) , (regs_regs_3_lpi_2[67:66])
      , (regs_regs_3_lpi_2[69:68]) , (regs_regs_3_lpi_2[71:70]) , (regs_regs_3_lpi_2[73:72])
      , (regs_regs_3_lpi_2[75:74]) , (regs_regs_3_lpi_2[77:76]) , (regs_regs_3_lpi_2[79:78])
      , (regs_regs_3_lpi_2[81:80]) , (regs_regs_3_lpi_2[83:82]) , (regs_regs_3_lpi_2[85:84])
      , (regs_regs_3_lpi_2[87:86]) , (regs_regs_3_lpi_2[89:88]) , (regs_regs_3_lpi_2[91:90])
      , (regs_regs_3_lpi_2[93:92]) , (regs_regs_3_lpi_2[95:94]) , (regs_regs_3_lpi_2[97:96])
      , (regs_regs_3_lpi_2[99:98]) , (regs_regs_3_lpi_2[101:100]) , (regs_regs_3_lpi_2[103:102])
      , (regs_regs_3_lpi_2[105:104]) , (regs_regs_3_lpi_2[107:106]) , (regs_regs_3_lpi_2[109:108])
      , (regs_regs_3_lpi_2[111:110]) , (regs_regs_3_lpi_2[113:112]) , (regs_regs_3_lpi_2[115:114])
      , (regs_regs_3_lpi_2[117:116]) , (regs_regs_3_lpi_2[119:118]) , (regs_regs_3_lpi_2[121:120])
      , (regs_regs_3_lpi_2[123:122]) , (regs_regs_3_lpi_2[125:124]) , (regs_regs_3_lpi_2[127:126])
      , (regs_regs_3_lpi_2[129:128]) , (regs_regs_3_lpi_2[131:130]) , (regs_regs_3_lpi_2[133:132])
      , (regs_regs_3_lpi_2[135:134]) , (regs_regs_3_lpi_2[137:136]) , (regs_regs_3_lpi_2[139:138])
      , (regs_regs_3_lpi_2[141:140]) , (regs_regs_3_lpi_2[143:142]) , (regs_regs_3_lpi_2[145:144])
      , (regs_regs_3_lpi_2[147:146]) , (regs_regs_3_lpi_2[149:148]) , (regs_regs_4_lpi_2[1:0])
      , (regs_regs_4_lpi_2[3:2]) , (regs_regs_4_lpi_2[5:4]) , (regs_regs_4_lpi_2[7:6])
      , (regs_regs_4_lpi_2[9:8]) , (regs_regs_4_lpi_2[11:10]) , (regs_regs_4_lpi_2[13:12])
      , (regs_regs_4_lpi_2[15:14]) , (regs_regs_4_lpi_2[17:16]) , (regs_regs_4_lpi_2[19:18])
      , (regs_regs_4_lpi_2[21:20]) , (regs_regs_4_lpi_2[23:22]) , (regs_regs_4_lpi_2[25:24])
      , (regs_regs_4_lpi_2[27:26]) , (regs_regs_4_lpi_2[29:28]) , (regs_regs_4_lpi_2[31:30])
      , (regs_regs_4_lpi_2[33:32]) , (regs_regs_4_lpi_2[35:34]) , (regs_regs_4_lpi_2[37:36])
      , (regs_regs_4_lpi_2[39:38]) , (regs_regs_4_lpi_2[41:40]) , (regs_regs_4_lpi_2[43:42])
      , (regs_regs_4_lpi_2[45:44]) , (regs_regs_4_lpi_2[47:46]) , (regs_regs_4_lpi_2[49:48])
      , (regs_regs_4_lpi_2[51:50]) , (regs_regs_4_lpi_2[53:52]) , (regs_regs_4_lpi_2[55:54])
      , (regs_regs_4_lpi_2[57:56]) , (regs_regs_4_lpi_2[59:58]) , (regs_regs_4_lpi_2[61:60])
      , (regs_regs_4_lpi_2[63:62]) , (regs_regs_4_lpi_2[65:64]) , (regs_regs_4_lpi_2[67:66])
      , (regs_regs_4_lpi_2[69:68]) , (regs_regs_4_lpi_2[71:70]) , (regs_regs_4_lpi_2[73:72])
      , (regs_regs_4_lpi_2[75:74]) , (regs_regs_4_lpi_2[77:76]) , (regs_regs_4_lpi_2[79:78])
      , (regs_regs_4_lpi_2[81:80]) , (regs_regs_4_lpi_2[83:82]) , (regs_regs_4_lpi_2[85:84])
      , (regs_regs_4_lpi_2[87:86]) , (regs_regs_4_lpi_2[89:88]) , (regs_regs_4_lpi_2[91:90])
      , (regs_regs_4_lpi_2[93:92]) , (regs_regs_4_lpi_2[95:94]) , (regs_regs_4_lpi_2[97:96])
      , (regs_regs_4_lpi_2[99:98]) , (regs_regs_4_lpi_2[101:100]) , (regs_regs_4_lpi_2[103:102])
      , (regs_regs_4_lpi_2[105:104]) , (regs_regs_4_lpi_2[107:106]) , (regs_regs_4_lpi_2[109:108])
      , (regs_regs_4_lpi_2[111:110]) , (regs_regs_4_lpi_2[113:112]) , (regs_regs_4_lpi_2[115:114])
      , (regs_regs_4_lpi_2[117:116]) , (regs_regs_4_lpi_2[119:118]) , (regs_regs_4_lpi_2[121:120])
      , (regs_regs_4_lpi_2[123:122]) , (regs_regs_4_lpi_2[125:124]) , (regs_regs_4_lpi_2[127:126])
      , (regs_regs_4_lpi_2[129:128]) , (regs_regs_4_lpi_2[131:130]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg4 = MUX_v_2_512_2({(regs_regs_0_lpi_2[9:8]) , (regs_regs_0_lpi_2[11:10])
      , (regs_regs_0_lpi_2[13:12]) , (regs_regs_0_lpi_2[15:14]) , (regs_regs_0_lpi_2[17:16])
      , (regs_regs_0_lpi_2[19:18]) , (regs_regs_0_lpi_2[21:20]) , (regs_regs_0_lpi_2[23:22])
      , (regs_regs_0_lpi_2[25:24]) , (regs_regs_0_lpi_2[27:26]) , (regs_regs_0_lpi_2[29:28])
      , (regs_regs_0_lpi_2[31:30]) , (regs_regs_0_lpi_2[33:32]) , (regs_regs_0_lpi_2[35:34])
      , (regs_regs_0_lpi_2[37:36]) , (regs_regs_0_lpi_2[39:38]) , (regs_regs_0_lpi_2[41:40])
      , (regs_regs_0_lpi_2[43:42]) , (regs_regs_0_lpi_2[45:44]) , (regs_regs_0_lpi_2[47:46])
      , (regs_regs_0_lpi_2[49:48]) , (regs_regs_0_lpi_2[51:50]) , (regs_regs_0_lpi_2[53:52])
      , (regs_regs_0_lpi_2[55:54]) , (regs_regs_0_lpi_2[57:56]) , (regs_regs_0_lpi_2[59:58])
      , (regs_regs_0_lpi_2[61:60]) , (regs_regs_0_lpi_2[63:62]) , (regs_regs_0_lpi_2[65:64])
      , (regs_regs_0_lpi_2[67:66]) , (regs_regs_0_lpi_2[69:68]) , (regs_regs_0_lpi_2[71:70])
      , (regs_regs_0_lpi_2[73:72]) , (regs_regs_0_lpi_2[75:74]) , (regs_regs_0_lpi_2[77:76])
      , (regs_regs_0_lpi_2[79:78]) , (regs_regs_0_lpi_2[81:80]) , (regs_regs_0_lpi_2[83:82])
      , (regs_regs_0_lpi_2[85:84]) , (regs_regs_0_lpi_2[87:86]) , (regs_regs_0_lpi_2[89:88])
      , (regs_regs_0_lpi_2[91:90]) , (regs_regs_0_lpi_2[93:92]) , (regs_regs_0_lpi_2[95:94])
      , (regs_regs_0_lpi_2[97:96]) , (regs_regs_0_lpi_2[99:98]) , (regs_regs_0_lpi_2[101:100])
      , (regs_regs_0_lpi_2[103:102]) , (regs_regs_0_lpi_2[105:104]) , (regs_regs_0_lpi_2[107:106])
      , (regs_regs_0_lpi_2[109:108]) , (regs_regs_0_lpi_2[111:110]) , (regs_regs_0_lpi_2[113:112])
      , (regs_regs_0_lpi_2[115:114]) , (regs_regs_0_lpi_2[117:116]) , (regs_regs_0_lpi_2[119:118])
      , (regs_regs_0_lpi_2[121:120]) , (regs_regs_0_lpi_2[123:122]) , (regs_regs_0_lpi_2[125:124])
      , (regs_regs_0_lpi_2[127:126]) , (regs_regs_0_lpi_2[129:128]) , (regs_regs_0_lpi_2[131:130])
      , (regs_regs_0_lpi_2[133:132]) , (regs_regs_0_lpi_2[135:134]) , (regs_regs_0_lpi_2[137:136])
      , (regs_regs_0_lpi_2[139:138]) , (regs_regs_0_lpi_2[141:140]) , (regs_regs_0_lpi_2[143:142])
      , (regs_regs_0_lpi_2[145:144]) , (regs_regs_0_lpi_2[147:146]) , (regs_regs_0_lpi_2[149:148])
      , (regs_regs_1_lpi_2[1:0]) , (regs_regs_1_lpi_2[3:2]) , (regs_regs_1_lpi_2[5:4])
      , (regs_regs_1_lpi_2[7:6]) , (regs_regs_1_lpi_2[9:8]) , (regs_regs_1_lpi_2[11:10])
      , (regs_regs_1_lpi_2[13:12]) , (regs_regs_1_lpi_2[15:14]) , (regs_regs_1_lpi_2[17:16])
      , (regs_regs_1_lpi_2[19:18]) , (regs_regs_1_lpi_2[21:20]) , (regs_regs_1_lpi_2[23:22])
      , (regs_regs_1_lpi_2[25:24]) , (regs_regs_1_lpi_2[27:26]) , (regs_regs_1_lpi_2[29:28])
      , (regs_regs_1_lpi_2[31:30]) , (regs_regs_1_lpi_2[33:32]) , (regs_regs_1_lpi_2[35:34])
      , (regs_regs_1_lpi_2[37:36]) , (regs_regs_1_lpi_2[39:38]) , (regs_regs_1_lpi_2[41:40])
      , (regs_regs_1_lpi_2[43:42]) , (regs_regs_1_lpi_2[45:44]) , (regs_regs_1_lpi_2[47:46])
      , (regs_regs_1_lpi_2[49:48]) , (regs_regs_1_lpi_2[51:50]) , (regs_regs_1_lpi_2[53:52])
      , (regs_regs_1_lpi_2[55:54]) , (regs_regs_1_lpi_2[57:56]) , (regs_regs_1_lpi_2[59:58])
      , (regs_regs_1_lpi_2[61:60]) , (regs_regs_1_lpi_2[63:62]) , (regs_regs_1_lpi_2[65:64])
      , (regs_regs_1_lpi_2[67:66]) , (regs_regs_1_lpi_2[69:68]) , (regs_regs_1_lpi_2[71:70])
      , (regs_regs_1_lpi_2[73:72]) , (regs_regs_1_lpi_2[75:74]) , (regs_regs_1_lpi_2[77:76])
      , (regs_regs_1_lpi_2[79:78]) , (regs_regs_1_lpi_2[81:80]) , (regs_regs_1_lpi_2[83:82])
      , (regs_regs_1_lpi_2[85:84]) , (regs_regs_1_lpi_2[87:86]) , (regs_regs_1_lpi_2[89:88])
      , (regs_regs_1_lpi_2[91:90]) , (regs_regs_1_lpi_2[93:92]) , (regs_regs_1_lpi_2[95:94])
      , (regs_regs_1_lpi_2[97:96]) , (regs_regs_1_lpi_2[99:98]) , (regs_regs_1_lpi_2[101:100])
      , (regs_regs_1_lpi_2[103:102]) , (regs_regs_1_lpi_2[105:104]) , (regs_regs_1_lpi_2[107:106])
      , (regs_regs_1_lpi_2[109:108]) , (regs_regs_1_lpi_2[111:110]) , (regs_regs_1_lpi_2[113:112])
      , (regs_regs_1_lpi_2[115:114]) , (regs_regs_1_lpi_2[117:116]) , (regs_regs_1_lpi_2[119:118])
      , (regs_regs_1_lpi_2[121:120]) , (regs_regs_1_lpi_2[123:122]) , (regs_regs_1_lpi_2[125:124])
      , (regs_regs_1_lpi_2[127:126]) , (regs_regs_1_lpi_2[129:128]) , (regs_regs_1_lpi_2[131:130])
      , (regs_regs_1_lpi_2[133:132]) , (regs_regs_1_lpi_2[135:134]) , (regs_regs_1_lpi_2[137:136])
      , (regs_regs_1_lpi_2[139:138]) , (regs_regs_1_lpi_2[141:140]) , (regs_regs_1_lpi_2[143:142])
      , (regs_regs_1_lpi_2[145:144]) , (regs_regs_1_lpi_2[147:146]) , (regs_regs_1_lpi_2[149:148])
      , (regs_regs_2_lpi_2[1:0]) , (regs_regs_2_lpi_2[3:2]) , (regs_regs_2_lpi_2[5:4])
      , (regs_regs_2_lpi_2[7:6]) , (regs_regs_2_lpi_2[9:8]) , (regs_regs_2_lpi_2[11:10])
      , (regs_regs_2_lpi_2[13:12]) , (regs_regs_2_lpi_2[15:14]) , (regs_regs_2_lpi_2[17:16])
      , (regs_regs_2_lpi_2[19:18]) , (regs_regs_2_lpi_2[21:20]) , (regs_regs_2_lpi_2[23:22])
      , (regs_regs_2_lpi_2[25:24]) , (regs_regs_2_lpi_2[27:26]) , (regs_regs_2_lpi_2[29:28])
      , (regs_regs_2_lpi_2[31:30]) , (regs_regs_2_lpi_2[33:32]) , (regs_regs_2_lpi_2[35:34])
      , (regs_regs_2_lpi_2[37:36]) , (regs_regs_2_lpi_2[39:38]) , (regs_regs_2_lpi_2[41:40])
      , (regs_regs_2_lpi_2[43:42]) , (regs_regs_2_lpi_2[45:44]) , (regs_regs_2_lpi_2[47:46])
      , (regs_regs_2_lpi_2[49:48]) , (regs_regs_2_lpi_2[51:50]) , (regs_regs_2_lpi_2[53:52])
      , (regs_regs_2_lpi_2[55:54]) , (regs_regs_2_lpi_2[57:56]) , (regs_regs_2_lpi_2[59:58])
      , (regs_regs_2_lpi_2[61:60]) , (regs_regs_2_lpi_2[63:62]) , (regs_regs_2_lpi_2[65:64])
      , (regs_regs_2_lpi_2[67:66]) , (regs_regs_2_lpi_2[69:68]) , (regs_regs_2_lpi_2[71:70])
      , (regs_regs_2_lpi_2[73:72]) , (regs_regs_2_lpi_2[75:74]) , (regs_regs_2_lpi_2[77:76])
      , (regs_regs_2_lpi_2[79:78]) , (regs_regs_2_lpi_2[81:80]) , (regs_regs_2_lpi_2[83:82])
      , (regs_regs_2_lpi_2[85:84]) , (regs_regs_2_lpi_2[87:86]) , (regs_regs_2_lpi_2[89:88])
      , (regs_regs_2_lpi_2[91:90]) , (regs_regs_2_lpi_2[93:92]) , (regs_regs_2_lpi_2[95:94])
      , (regs_regs_2_lpi_2[97:96]) , (regs_regs_2_lpi_2[99:98]) , (regs_regs_2_lpi_2[101:100])
      , (regs_regs_2_lpi_2[103:102]) , (regs_regs_2_lpi_2[105:104]) , (regs_regs_2_lpi_2[107:106])
      , (regs_regs_2_lpi_2[109:108]) , (regs_regs_2_lpi_2[111:110]) , (regs_regs_2_lpi_2[113:112])
      , (regs_regs_2_lpi_2[115:114]) , (regs_regs_2_lpi_2[117:116]) , (regs_regs_2_lpi_2[119:118])
      , (regs_regs_2_lpi_2[121:120]) , (regs_regs_2_lpi_2[123:122]) , (regs_regs_2_lpi_2[125:124])
      , (regs_regs_2_lpi_2[127:126]) , (regs_regs_2_lpi_2[129:128]) , (regs_regs_2_lpi_2[131:130])
      , (regs_regs_2_lpi_2[133:132]) , (regs_regs_2_lpi_2[135:134]) , (regs_regs_2_lpi_2[137:136])
      , (regs_regs_2_lpi_2[139:138]) , (regs_regs_2_lpi_2[141:140]) , (regs_regs_2_lpi_2[143:142])
      , (regs_regs_2_lpi_2[145:144]) , (regs_regs_2_lpi_2[147:146]) , (regs_regs_2_lpi_2[149:148])
      , (regs_regs_3_lpi_2[1:0]) , (regs_regs_3_lpi_2[3:2]) , (regs_regs_3_lpi_2[5:4])
      , (regs_regs_3_lpi_2[7:6]) , (regs_regs_3_lpi_2[9:8]) , (regs_regs_3_lpi_2[11:10])
      , (regs_regs_3_lpi_2[13:12]) , (regs_regs_3_lpi_2[15:14]) , (regs_regs_3_lpi_2[17:16])
      , (regs_regs_3_lpi_2[19:18]) , (regs_regs_3_lpi_2[21:20]) , (regs_regs_3_lpi_2[23:22])
      , (regs_regs_3_lpi_2[25:24]) , (regs_regs_3_lpi_2[27:26]) , (regs_regs_3_lpi_2[29:28])
      , (regs_regs_3_lpi_2[31:30]) , (regs_regs_3_lpi_2[33:32]) , (regs_regs_3_lpi_2[35:34])
      , (regs_regs_3_lpi_2[37:36]) , (regs_regs_3_lpi_2[39:38]) , (regs_regs_3_lpi_2[41:40])
      , (regs_regs_3_lpi_2[43:42]) , (regs_regs_3_lpi_2[45:44]) , (regs_regs_3_lpi_2[47:46])
      , (regs_regs_3_lpi_2[49:48]) , (regs_regs_3_lpi_2[51:50]) , (regs_regs_3_lpi_2[53:52])
      , (regs_regs_3_lpi_2[55:54]) , (regs_regs_3_lpi_2[57:56]) , (regs_regs_3_lpi_2[59:58])
      , (regs_regs_3_lpi_2[61:60]) , (regs_regs_3_lpi_2[63:62]) , (regs_regs_3_lpi_2[65:64])
      , (regs_regs_3_lpi_2[67:66]) , (regs_regs_3_lpi_2[69:68]) , (regs_regs_3_lpi_2[71:70])
      , (regs_regs_3_lpi_2[73:72]) , (regs_regs_3_lpi_2[75:74]) , (regs_regs_3_lpi_2[77:76])
      , (regs_regs_3_lpi_2[79:78]) , (regs_regs_3_lpi_2[81:80]) , (regs_regs_3_lpi_2[83:82])
      , (regs_regs_3_lpi_2[85:84]) , (regs_regs_3_lpi_2[87:86]) , (regs_regs_3_lpi_2[89:88])
      , (regs_regs_3_lpi_2[91:90]) , (regs_regs_3_lpi_2[93:92]) , (regs_regs_3_lpi_2[95:94])
      , (regs_regs_3_lpi_2[97:96]) , (regs_regs_3_lpi_2[99:98]) , (regs_regs_3_lpi_2[101:100])
      , (regs_regs_3_lpi_2[103:102]) , (regs_regs_3_lpi_2[105:104]) , (regs_regs_3_lpi_2[107:106])
      , (regs_regs_3_lpi_2[109:108]) , (regs_regs_3_lpi_2[111:110]) , (regs_regs_3_lpi_2[113:112])
      , (regs_regs_3_lpi_2[115:114]) , (regs_regs_3_lpi_2[117:116]) , (regs_regs_3_lpi_2[119:118])
      , (regs_regs_3_lpi_2[121:120]) , (regs_regs_3_lpi_2[123:122]) , (regs_regs_3_lpi_2[125:124])
      , (regs_regs_3_lpi_2[127:126]) , (regs_regs_3_lpi_2[129:128]) , (regs_regs_3_lpi_2[131:130])
      , (regs_regs_3_lpi_2[133:132]) , (regs_regs_3_lpi_2[135:134]) , (regs_regs_3_lpi_2[137:136])
      , (regs_regs_3_lpi_2[139:138]) , (regs_regs_3_lpi_2[141:140]) , (regs_regs_3_lpi_2[143:142])
      , (regs_regs_3_lpi_2[145:144]) , (regs_regs_3_lpi_2[147:146]) , (regs_regs_3_lpi_2[149:148])
      , (regs_regs_4_lpi_2[1:0]) , (regs_regs_4_lpi_2[3:2]) , (regs_regs_4_lpi_2[5:4])
      , (regs_regs_4_lpi_2[7:6]) , (regs_regs_4_lpi_2[9:8]) , (regs_regs_4_lpi_2[11:10])
      , (regs_regs_4_lpi_2[13:12]) , (regs_regs_4_lpi_2[15:14]) , (regs_regs_4_lpi_2[17:16])
      , (regs_regs_4_lpi_2[19:18]) , (regs_regs_4_lpi_2[21:20]) , (regs_regs_4_lpi_2[23:22])
      , (regs_regs_4_lpi_2[25:24]) , (regs_regs_4_lpi_2[27:26]) , (regs_regs_4_lpi_2[29:28])
      , (regs_regs_4_lpi_2[31:30]) , (regs_regs_4_lpi_2[33:32]) , (regs_regs_4_lpi_2[35:34])
      , (regs_regs_4_lpi_2[37:36]) , (regs_regs_4_lpi_2[39:38]) , (regs_regs_4_lpi_2[41:40])
      , (regs_regs_4_lpi_2[43:42]) , (regs_regs_4_lpi_2[45:44]) , (regs_regs_4_lpi_2[47:46])
      , (regs_regs_4_lpi_2[49:48]) , (regs_regs_4_lpi_2[51:50]) , (regs_regs_4_lpi_2[53:52])
      , (regs_regs_4_lpi_2[55:54]) , (regs_regs_4_lpi_2[57:56]) , (regs_regs_4_lpi_2[59:58])
      , (regs_regs_4_lpi_2[61:60]) , (regs_regs_4_lpi_2[63:62]) , (regs_regs_4_lpi_2[65:64])
      , (regs_regs_4_lpi_2[67:66]) , (regs_regs_4_lpi_2[69:68]) , (regs_regs_4_lpi_2[71:70])
      , (regs_regs_4_lpi_2[73:72]) , (regs_regs_4_lpi_2[75:74]) , (regs_regs_4_lpi_2[77:76])
      , (regs_regs_4_lpi_2[79:78]) , (regs_regs_4_lpi_2[81:80]) , (regs_regs_4_lpi_2[83:82])
      , (regs_regs_4_lpi_2[85:84]) , (regs_regs_4_lpi_2[87:86]) , (regs_regs_4_lpi_2[89:88])
      , (regs_regs_4_lpi_2[91:90]) , (regs_regs_4_lpi_2[93:92]) , (regs_regs_4_lpi_2[95:94])
      , (regs_regs_4_lpi_2[97:96]) , (regs_regs_4_lpi_2[99:98]) , (regs_regs_4_lpi_2[101:100])
      , (regs_regs_4_lpi_2[103:102]) , (regs_regs_4_lpi_2[105:104]) , (regs_regs_4_lpi_2[107:106])
      , (regs_regs_4_lpi_2[109:108]) , (regs_regs_4_lpi_2[111:110]) , (regs_regs_4_lpi_2[113:112])
      , (regs_regs_4_lpi_2[115:114]) , (regs_regs_4_lpi_2[117:116]) , (regs_regs_4_lpi_2[119:118])
      , (regs_regs_4_lpi_2[121:120]) , (regs_regs_4_lpi_2[123:122]) , (regs_regs_4_lpi_2[125:124])
      , (regs_regs_4_lpi_2[127:126]) , (regs_regs_4_lpi_2[129:128]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg3 = MUX_v_2_512_2({(regs_regs_0_lpi_2[7:6]) , (regs_regs_0_lpi_2[9:8])
      , (regs_regs_0_lpi_2[11:10]) , (regs_regs_0_lpi_2[13:12]) , (regs_regs_0_lpi_2[15:14])
      , (regs_regs_0_lpi_2[17:16]) , (regs_regs_0_lpi_2[19:18]) , (regs_regs_0_lpi_2[21:20])
      , (regs_regs_0_lpi_2[23:22]) , (regs_regs_0_lpi_2[25:24]) , (regs_regs_0_lpi_2[27:26])
      , (regs_regs_0_lpi_2[29:28]) , (regs_regs_0_lpi_2[31:30]) , (regs_regs_0_lpi_2[33:32])
      , (regs_regs_0_lpi_2[35:34]) , (regs_regs_0_lpi_2[37:36]) , (regs_regs_0_lpi_2[39:38])
      , (regs_regs_0_lpi_2[41:40]) , (regs_regs_0_lpi_2[43:42]) , (regs_regs_0_lpi_2[45:44])
      , (regs_regs_0_lpi_2[47:46]) , (regs_regs_0_lpi_2[49:48]) , (regs_regs_0_lpi_2[51:50])
      , (regs_regs_0_lpi_2[53:52]) , (regs_regs_0_lpi_2[55:54]) , (regs_regs_0_lpi_2[57:56])
      , (regs_regs_0_lpi_2[59:58]) , (regs_regs_0_lpi_2[61:60]) , (regs_regs_0_lpi_2[63:62])
      , (regs_regs_0_lpi_2[65:64]) , (regs_regs_0_lpi_2[67:66]) , (regs_regs_0_lpi_2[69:68])
      , (regs_regs_0_lpi_2[71:70]) , (regs_regs_0_lpi_2[73:72]) , (regs_regs_0_lpi_2[75:74])
      , (regs_regs_0_lpi_2[77:76]) , (regs_regs_0_lpi_2[79:78]) , (regs_regs_0_lpi_2[81:80])
      , (regs_regs_0_lpi_2[83:82]) , (regs_regs_0_lpi_2[85:84]) , (regs_regs_0_lpi_2[87:86])
      , (regs_regs_0_lpi_2[89:88]) , (regs_regs_0_lpi_2[91:90]) , (regs_regs_0_lpi_2[93:92])
      , (regs_regs_0_lpi_2[95:94]) , (regs_regs_0_lpi_2[97:96]) , (regs_regs_0_lpi_2[99:98])
      , (regs_regs_0_lpi_2[101:100]) , (regs_regs_0_lpi_2[103:102]) , (regs_regs_0_lpi_2[105:104])
      , (regs_regs_0_lpi_2[107:106]) , (regs_regs_0_lpi_2[109:108]) , (regs_regs_0_lpi_2[111:110])
      , (regs_regs_0_lpi_2[113:112]) , (regs_regs_0_lpi_2[115:114]) , (regs_regs_0_lpi_2[117:116])
      , (regs_regs_0_lpi_2[119:118]) , (regs_regs_0_lpi_2[121:120]) , (regs_regs_0_lpi_2[123:122])
      , (regs_regs_0_lpi_2[125:124]) , (regs_regs_0_lpi_2[127:126]) , (regs_regs_0_lpi_2[129:128])
      , (regs_regs_0_lpi_2[131:130]) , (regs_regs_0_lpi_2[133:132]) , (regs_regs_0_lpi_2[135:134])
      , (regs_regs_0_lpi_2[137:136]) , (regs_regs_0_lpi_2[139:138]) , (regs_regs_0_lpi_2[141:140])
      , (regs_regs_0_lpi_2[143:142]) , (regs_regs_0_lpi_2[145:144]) , (regs_regs_0_lpi_2[147:146])
      , (regs_regs_0_lpi_2[149:148]) , (regs_regs_1_lpi_2[1:0]) , (regs_regs_1_lpi_2[3:2])
      , (regs_regs_1_lpi_2[5:4]) , (regs_regs_1_lpi_2[7:6]) , (regs_regs_1_lpi_2[9:8])
      , (regs_regs_1_lpi_2[11:10]) , (regs_regs_1_lpi_2[13:12]) , (regs_regs_1_lpi_2[15:14])
      , (regs_regs_1_lpi_2[17:16]) , (regs_regs_1_lpi_2[19:18]) , (regs_regs_1_lpi_2[21:20])
      , (regs_regs_1_lpi_2[23:22]) , (regs_regs_1_lpi_2[25:24]) , (regs_regs_1_lpi_2[27:26])
      , (regs_regs_1_lpi_2[29:28]) , (regs_regs_1_lpi_2[31:30]) , (regs_regs_1_lpi_2[33:32])
      , (regs_regs_1_lpi_2[35:34]) , (regs_regs_1_lpi_2[37:36]) , (regs_regs_1_lpi_2[39:38])
      , (regs_regs_1_lpi_2[41:40]) , (regs_regs_1_lpi_2[43:42]) , (regs_regs_1_lpi_2[45:44])
      , (regs_regs_1_lpi_2[47:46]) , (regs_regs_1_lpi_2[49:48]) , (regs_regs_1_lpi_2[51:50])
      , (regs_regs_1_lpi_2[53:52]) , (regs_regs_1_lpi_2[55:54]) , (regs_regs_1_lpi_2[57:56])
      , (regs_regs_1_lpi_2[59:58]) , (regs_regs_1_lpi_2[61:60]) , (regs_regs_1_lpi_2[63:62])
      , (regs_regs_1_lpi_2[65:64]) , (regs_regs_1_lpi_2[67:66]) , (regs_regs_1_lpi_2[69:68])
      , (regs_regs_1_lpi_2[71:70]) , (regs_regs_1_lpi_2[73:72]) , (regs_regs_1_lpi_2[75:74])
      , (regs_regs_1_lpi_2[77:76]) , (regs_regs_1_lpi_2[79:78]) , (regs_regs_1_lpi_2[81:80])
      , (regs_regs_1_lpi_2[83:82]) , (regs_regs_1_lpi_2[85:84]) , (regs_regs_1_lpi_2[87:86])
      , (regs_regs_1_lpi_2[89:88]) , (regs_regs_1_lpi_2[91:90]) , (regs_regs_1_lpi_2[93:92])
      , (regs_regs_1_lpi_2[95:94]) , (regs_regs_1_lpi_2[97:96]) , (regs_regs_1_lpi_2[99:98])
      , (regs_regs_1_lpi_2[101:100]) , (regs_regs_1_lpi_2[103:102]) , (regs_regs_1_lpi_2[105:104])
      , (regs_regs_1_lpi_2[107:106]) , (regs_regs_1_lpi_2[109:108]) , (regs_regs_1_lpi_2[111:110])
      , (regs_regs_1_lpi_2[113:112]) , (regs_regs_1_lpi_2[115:114]) , (regs_regs_1_lpi_2[117:116])
      , (regs_regs_1_lpi_2[119:118]) , (regs_regs_1_lpi_2[121:120]) , (regs_regs_1_lpi_2[123:122])
      , (regs_regs_1_lpi_2[125:124]) , (regs_regs_1_lpi_2[127:126]) , (regs_regs_1_lpi_2[129:128])
      , (regs_regs_1_lpi_2[131:130]) , (regs_regs_1_lpi_2[133:132]) , (regs_regs_1_lpi_2[135:134])
      , (regs_regs_1_lpi_2[137:136]) , (regs_regs_1_lpi_2[139:138]) , (regs_regs_1_lpi_2[141:140])
      , (regs_regs_1_lpi_2[143:142]) , (regs_regs_1_lpi_2[145:144]) , (regs_regs_1_lpi_2[147:146])
      , (regs_regs_1_lpi_2[149:148]) , (regs_regs_2_lpi_2[1:0]) , (regs_regs_2_lpi_2[3:2])
      , (regs_regs_2_lpi_2[5:4]) , (regs_regs_2_lpi_2[7:6]) , (regs_regs_2_lpi_2[9:8])
      , (regs_regs_2_lpi_2[11:10]) , (regs_regs_2_lpi_2[13:12]) , (regs_regs_2_lpi_2[15:14])
      , (regs_regs_2_lpi_2[17:16]) , (regs_regs_2_lpi_2[19:18]) , (regs_regs_2_lpi_2[21:20])
      , (regs_regs_2_lpi_2[23:22]) , (regs_regs_2_lpi_2[25:24]) , (regs_regs_2_lpi_2[27:26])
      , (regs_regs_2_lpi_2[29:28]) , (regs_regs_2_lpi_2[31:30]) , (regs_regs_2_lpi_2[33:32])
      , (regs_regs_2_lpi_2[35:34]) , (regs_regs_2_lpi_2[37:36]) , (regs_regs_2_lpi_2[39:38])
      , (regs_regs_2_lpi_2[41:40]) , (regs_regs_2_lpi_2[43:42]) , (regs_regs_2_lpi_2[45:44])
      , (regs_regs_2_lpi_2[47:46]) , (regs_regs_2_lpi_2[49:48]) , (regs_regs_2_lpi_2[51:50])
      , (regs_regs_2_lpi_2[53:52]) , (regs_regs_2_lpi_2[55:54]) , (regs_regs_2_lpi_2[57:56])
      , (regs_regs_2_lpi_2[59:58]) , (regs_regs_2_lpi_2[61:60]) , (regs_regs_2_lpi_2[63:62])
      , (regs_regs_2_lpi_2[65:64]) , (regs_regs_2_lpi_2[67:66]) , (regs_regs_2_lpi_2[69:68])
      , (regs_regs_2_lpi_2[71:70]) , (regs_regs_2_lpi_2[73:72]) , (regs_regs_2_lpi_2[75:74])
      , (regs_regs_2_lpi_2[77:76]) , (regs_regs_2_lpi_2[79:78]) , (regs_regs_2_lpi_2[81:80])
      , (regs_regs_2_lpi_2[83:82]) , (regs_regs_2_lpi_2[85:84]) , (regs_regs_2_lpi_2[87:86])
      , (regs_regs_2_lpi_2[89:88]) , (regs_regs_2_lpi_2[91:90]) , (regs_regs_2_lpi_2[93:92])
      , (regs_regs_2_lpi_2[95:94]) , (regs_regs_2_lpi_2[97:96]) , (regs_regs_2_lpi_2[99:98])
      , (regs_regs_2_lpi_2[101:100]) , (regs_regs_2_lpi_2[103:102]) , (regs_regs_2_lpi_2[105:104])
      , (regs_regs_2_lpi_2[107:106]) , (regs_regs_2_lpi_2[109:108]) , (regs_regs_2_lpi_2[111:110])
      , (regs_regs_2_lpi_2[113:112]) , (regs_regs_2_lpi_2[115:114]) , (regs_regs_2_lpi_2[117:116])
      , (regs_regs_2_lpi_2[119:118]) , (regs_regs_2_lpi_2[121:120]) , (regs_regs_2_lpi_2[123:122])
      , (regs_regs_2_lpi_2[125:124]) , (regs_regs_2_lpi_2[127:126]) , (regs_regs_2_lpi_2[129:128])
      , (regs_regs_2_lpi_2[131:130]) , (regs_regs_2_lpi_2[133:132]) , (regs_regs_2_lpi_2[135:134])
      , (regs_regs_2_lpi_2[137:136]) , (regs_regs_2_lpi_2[139:138]) , (regs_regs_2_lpi_2[141:140])
      , (regs_regs_2_lpi_2[143:142]) , (regs_regs_2_lpi_2[145:144]) , (regs_regs_2_lpi_2[147:146])
      , (regs_regs_2_lpi_2[149:148]) , (regs_regs_3_lpi_2[1:0]) , (regs_regs_3_lpi_2[3:2])
      , (regs_regs_3_lpi_2[5:4]) , (regs_regs_3_lpi_2[7:6]) , (regs_regs_3_lpi_2[9:8])
      , (regs_regs_3_lpi_2[11:10]) , (regs_regs_3_lpi_2[13:12]) , (regs_regs_3_lpi_2[15:14])
      , (regs_regs_3_lpi_2[17:16]) , (regs_regs_3_lpi_2[19:18]) , (regs_regs_3_lpi_2[21:20])
      , (regs_regs_3_lpi_2[23:22]) , (regs_regs_3_lpi_2[25:24]) , (regs_regs_3_lpi_2[27:26])
      , (regs_regs_3_lpi_2[29:28]) , (regs_regs_3_lpi_2[31:30]) , (regs_regs_3_lpi_2[33:32])
      , (regs_regs_3_lpi_2[35:34]) , (regs_regs_3_lpi_2[37:36]) , (regs_regs_3_lpi_2[39:38])
      , (regs_regs_3_lpi_2[41:40]) , (regs_regs_3_lpi_2[43:42]) , (regs_regs_3_lpi_2[45:44])
      , (regs_regs_3_lpi_2[47:46]) , (regs_regs_3_lpi_2[49:48]) , (regs_regs_3_lpi_2[51:50])
      , (regs_regs_3_lpi_2[53:52]) , (regs_regs_3_lpi_2[55:54]) , (regs_regs_3_lpi_2[57:56])
      , (regs_regs_3_lpi_2[59:58]) , (regs_regs_3_lpi_2[61:60]) , (regs_regs_3_lpi_2[63:62])
      , (regs_regs_3_lpi_2[65:64]) , (regs_regs_3_lpi_2[67:66]) , (regs_regs_3_lpi_2[69:68])
      , (regs_regs_3_lpi_2[71:70]) , (regs_regs_3_lpi_2[73:72]) , (regs_regs_3_lpi_2[75:74])
      , (regs_regs_3_lpi_2[77:76]) , (regs_regs_3_lpi_2[79:78]) , (regs_regs_3_lpi_2[81:80])
      , (regs_regs_3_lpi_2[83:82]) , (regs_regs_3_lpi_2[85:84]) , (regs_regs_3_lpi_2[87:86])
      , (regs_regs_3_lpi_2[89:88]) , (regs_regs_3_lpi_2[91:90]) , (regs_regs_3_lpi_2[93:92])
      , (regs_regs_3_lpi_2[95:94]) , (regs_regs_3_lpi_2[97:96]) , (regs_regs_3_lpi_2[99:98])
      , (regs_regs_3_lpi_2[101:100]) , (regs_regs_3_lpi_2[103:102]) , (regs_regs_3_lpi_2[105:104])
      , (regs_regs_3_lpi_2[107:106]) , (regs_regs_3_lpi_2[109:108]) , (regs_regs_3_lpi_2[111:110])
      , (regs_regs_3_lpi_2[113:112]) , (regs_regs_3_lpi_2[115:114]) , (regs_regs_3_lpi_2[117:116])
      , (regs_regs_3_lpi_2[119:118]) , (regs_regs_3_lpi_2[121:120]) , (regs_regs_3_lpi_2[123:122])
      , (regs_regs_3_lpi_2[125:124]) , (regs_regs_3_lpi_2[127:126]) , (regs_regs_3_lpi_2[129:128])
      , (regs_regs_3_lpi_2[131:130]) , (regs_regs_3_lpi_2[133:132]) , (regs_regs_3_lpi_2[135:134])
      , (regs_regs_3_lpi_2[137:136]) , (regs_regs_3_lpi_2[139:138]) , (regs_regs_3_lpi_2[141:140])
      , (regs_regs_3_lpi_2[143:142]) , (regs_regs_3_lpi_2[145:144]) , (regs_regs_3_lpi_2[147:146])
      , (regs_regs_3_lpi_2[149:148]) , (regs_regs_4_lpi_2[1:0]) , (regs_regs_4_lpi_2[3:2])
      , (regs_regs_4_lpi_2[5:4]) , (regs_regs_4_lpi_2[7:6]) , (regs_regs_4_lpi_2[9:8])
      , (regs_regs_4_lpi_2[11:10]) , (regs_regs_4_lpi_2[13:12]) , (regs_regs_4_lpi_2[15:14])
      , (regs_regs_4_lpi_2[17:16]) , (regs_regs_4_lpi_2[19:18]) , (regs_regs_4_lpi_2[21:20])
      , (regs_regs_4_lpi_2[23:22]) , (regs_regs_4_lpi_2[25:24]) , (regs_regs_4_lpi_2[27:26])
      , (regs_regs_4_lpi_2[29:28]) , (regs_regs_4_lpi_2[31:30]) , (regs_regs_4_lpi_2[33:32])
      , (regs_regs_4_lpi_2[35:34]) , (regs_regs_4_lpi_2[37:36]) , (regs_regs_4_lpi_2[39:38])
      , (regs_regs_4_lpi_2[41:40]) , (regs_regs_4_lpi_2[43:42]) , (regs_regs_4_lpi_2[45:44])
      , (regs_regs_4_lpi_2[47:46]) , (regs_regs_4_lpi_2[49:48]) , (regs_regs_4_lpi_2[51:50])
      , (regs_regs_4_lpi_2[53:52]) , (regs_regs_4_lpi_2[55:54]) , (regs_regs_4_lpi_2[57:56])
      , (regs_regs_4_lpi_2[59:58]) , (regs_regs_4_lpi_2[61:60]) , (regs_regs_4_lpi_2[63:62])
      , (regs_regs_4_lpi_2[65:64]) , (regs_regs_4_lpi_2[67:66]) , (regs_regs_4_lpi_2[69:68])
      , (regs_regs_4_lpi_2[71:70]) , (regs_regs_4_lpi_2[73:72]) , (regs_regs_4_lpi_2[75:74])
      , (regs_regs_4_lpi_2[77:76]) , (regs_regs_4_lpi_2[79:78]) , (regs_regs_4_lpi_2[81:80])
      , (regs_regs_4_lpi_2[83:82]) , (regs_regs_4_lpi_2[85:84]) , (regs_regs_4_lpi_2[87:86])
      , (regs_regs_4_lpi_2[89:88]) , (regs_regs_4_lpi_2[91:90]) , (regs_regs_4_lpi_2[93:92])
      , (regs_regs_4_lpi_2[95:94]) , (regs_regs_4_lpi_2[97:96]) , (regs_regs_4_lpi_2[99:98])
      , (regs_regs_4_lpi_2[101:100]) , (regs_regs_4_lpi_2[103:102]) , (regs_regs_4_lpi_2[105:104])
      , (regs_regs_4_lpi_2[107:106]) , (regs_regs_4_lpi_2[109:108]) , (regs_regs_4_lpi_2[111:110])
      , (regs_regs_4_lpi_2[113:112]) , (regs_regs_4_lpi_2[115:114]) , (regs_regs_4_lpi_2[117:116])
      , (regs_regs_4_lpi_2[119:118]) , (regs_regs_4_lpi_2[121:120]) , (regs_regs_4_lpi_2[123:122])
      , (regs_regs_4_lpi_2[125:124]) , (regs_regs_4_lpi_2[127:126]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg2 = MUX_v_2_512_2({(regs_regs_0_lpi_2[5:4]) , (regs_regs_0_lpi_2[7:6])
      , (regs_regs_0_lpi_2[9:8]) , (regs_regs_0_lpi_2[11:10]) , (regs_regs_0_lpi_2[13:12])
      , (regs_regs_0_lpi_2[15:14]) , (regs_regs_0_lpi_2[17:16]) , (regs_regs_0_lpi_2[19:18])
      , (regs_regs_0_lpi_2[21:20]) , (regs_regs_0_lpi_2[23:22]) , (regs_regs_0_lpi_2[25:24])
      , (regs_regs_0_lpi_2[27:26]) , (regs_regs_0_lpi_2[29:28]) , (regs_regs_0_lpi_2[31:30])
      , (regs_regs_0_lpi_2[33:32]) , (regs_regs_0_lpi_2[35:34]) , (regs_regs_0_lpi_2[37:36])
      , (regs_regs_0_lpi_2[39:38]) , (regs_regs_0_lpi_2[41:40]) , (regs_regs_0_lpi_2[43:42])
      , (regs_regs_0_lpi_2[45:44]) , (regs_regs_0_lpi_2[47:46]) , (regs_regs_0_lpi_2[49:48])
      , (regs_regs_0_lpi_2[51:50]) , (regs_regs_0_lpi_2[53:52]) , (regs_regs_0_lpi_2[55:54])
      , (regs_regs_0_lpi_2[57:56]) , (regs_regs_0_lpi_2[59:58]) , (regs_regs_0_lpi_2[61:60])
      , (regs_regs_0_lpi_2[63:62]) , (regs_regs_0_lpi_2[65:64]) , (regs_regs_0_lpi_2[67:66])
      , (regs_regs_0_lpi_2[69:68]) , (regs_regs_0_lpi_2[71:70]) , (regs_regs_0_lpi_2[73:72])
      , (regs_regs_0_lpi_2[75:74]) , (regs_regs_0_lpi_2[77:76]) , (regs_regs_0_lpi_2[79:78])
      , (regs_regs_0_lpi_2[81:80]) , (regs_regs_0_lpi_2[83:82]) , (regs_regs_0_lpi_2[85:84])
      , (regs_regs_0_lpi_2[87:86]) , (regs_regs_0_lpi_2[89:88]) , (regs_regs_0_lpi_2[91:90])
      , (regs_regs_0_lpi_2[93:92]) , (regs_regs_0_lpi_2[95:94]) , (regs_regs_0_lpi_2[97:96])
      , (regs_regs_0_lpi_2[99:98]) , (regs_regs_0_lpi_2[101:100]) , (regs_regs_0_lpi_2[103:102])
      , (regs_regs_0_lpi_2[105:104]) , (regs_regs_0_lpi_2[107:106]) , (regs_regs_0_lpi_2[109:108])
      , (regs_regs_0_lpi_2[111:110]) , (regs_regs_0_lpi_2[113:112]) , (regs_regs_0_lpi_2[115:114])
      , (regs_regs_0_lpi_2[117:116]) , (regs_regs_0_lpi_2[119:118]) , (regs_regs_0_lpi_2[121:120])
      , (regs_regs_0_lpi_2[123:122]) , (regs_regs_0_lpi_2[125:124]) , (regs_regs_0_lpi_2[127:126])
      , (regs_regs_0_lpi_2[129:128]) , (regs_regs_0_lpi_2[131:130]) , (regs_regs_0_lpi_2[133:132])
      , (regs_regs_0_lpi_2[135:134]) , (regs_regs_0_lpi_2[137:136]) , (regs_regs_0_lpi_2[139:138])
      , (regs_regs_0_lpi_2[141:140]) , (regs_regs_0_lpi_2[143:142]) , (regs_regs_0_lpi_2[145:144])
      , (regs_regs_0_lpi_2[147:146]) , (regs_regs_0_lpi_2[149:148]) , (regs_regs_1_lpi_2[1:0])
      , (regs_regs_1_lpi_2[3:2]) , (regs_regs_1_lpi_2[5:4]) , (regs_regs_1_lpi_2[7:6])
      , (regs_regs_1_lpi_2[9:8]) , (regs_regs_1_lpi_2[11:10]) , (regs_regs_1_lpi_2[13:12])
      , (regs_regs_1_lpi_2[15:14]) , (regs_regs_1_lpi_2[17:16]) , (regs_regs_1_lpi_2[19:18])
      , (regs_regs_1_lpi_2[21:20]) , (regs_regs_1_lpi_2[23:22]) , (regs_regs_1_lpi_2[25:24])
      , (regs_regs_1_lpi_2[27:26]) , (regs_regs_1_lpi_2[29:28]) , (regs_regs_1_lpi_2[31:30])
      , (regs_regs_1_lpi_2[33:32]) , (regs_regs_1_lpi_2[35:34]) , (regs_regs_1_lpi_2[37:36])
      , (regs_regs_1_lpi_2[39:38]) , (regs_regs_1_lpi_2[41:40]) , (regs_regs_1_lpi_2[43:42])
      , (regs_regs_1_lpi_2[45:44]) , (regs_regs_1_lpi_2[47:46]) , (regs_regs_1_lpi_2[49:48])
      , (regs_regs_1_lpi_2[51:50]) , (regs_regs_1_lpi_2[53:52]) , (regs_regs_1_lpi_2[55:54])
      , (regs_regs_1_lpi_2[57:56]) , (regs_regs_1_lpi_2[59:58]) , (regs_regs_1_lpi_2[61:60])
      , (regs_regs_1_lpi_2[63:62]) , (regs_regs_1_lpi_2[65:64]) , (regs_regs_1_lpi_2[67:66])
      , (regs_regs_1_lpi_2[69:68]) , (regs_regs_1_lpi_2[71:70]) , (regs_regs_1_lpi_2[73:72])
      , (regs_regs_1_lpi_2[75:74]) , (regs_regs_1_lpi_2[77:76]) , (regs_regs_1_lpi_2[79:78])
      , (regs_regs_1_lpi_2[81:80]) , (regs_regs_1_lpi_2[83:82]) , (regs_regs_1_lpi_2[85:84])
      , (regs_regs_1_lpi_2[87:86]) , (regs_regs_1_lpi_2[89:88]) , (regs_regs_1_lpi_2[91:90])
      , (regs_regs_1_lpi_2[93:92]) , (regs_regs_1_lpi_2[95:94]) , (regs_regs_1_lpi_2[97:96])
      , (regs_regs_1_lpi_2[99:98]) , (regs_regs_1_lpi_2[101:100]) , (regs_regs_1_lpi_2[103:102])
      , (regs_regs_1_lpi_2[105:104]) , (regs_regs_1_lpi_2[107:106]) , (regs_regs_1_lpi_2[109:108])
      , (regs_regs_1_lpi_2[111:110]) , (regs_regs_1_lpi_2[113:112]) , (regs_regs_1_lpi_2[115:114])
      , (regs_regs_1_lpi_2[117:116]) , (regs_regs_1_lpi_2[119:118]) , (regs_regs_1_lpi_2[121:120])
      , (regs_regs_1_lpi_2[123:122]) , (regs_regs_1_lpi_2[125:124]) , (regs_regs_1_lpi_2[127:126])
      , (regs_regs_1_lpi_2[129:128]) , (regs_regs_1_lpi_2[131:130]) , (regs_regs_1_lpi_2[133:132])
      , (regs_regs_1_lpi_2[135:134]) , (regs_regs_1_lpi_2[137:136]) , (regs_regs_1_lpi_2[139:138])
      , (regs_regs_1_lpi_2[141:140]) , (regs_regs_1_lpi_2[143:142]) , (regs_regs_1_lpi_2[145:144])
      , (regs_regs_1_lpi_2[147:146]) , (regs_regs_1_lpi_2[149:148]) , (regs_regs_2_lpi_2[1:0])
      , (regs_regs_2_lpi_2[3:2]) , (regs_regs_2_lpi_2[5:4]) , (regs_regs_2_lpi_2[7:6])
      , (regs_regs_2_lpi_2[9:8]) , (regs_regs_2_lpi_2[11:10]) , (regs_regs_2_lpi_2[13:12])
      , (regs_regs_2_lpi_2[15:14]) , (regs_regs_2_lpi_2[17:16]) , (regs_regs_2_lpi_2[19:18])
      , (regs_regs_2_lpi_2[21:20]) , (regs_regs_2_lpi_2[23:22]) , (regs_regs_2_lpi_2[25:24])
      , (regs_regs_2_lpi_2[27:26]) , (regs_regs_2_lpi_2[29:28]) , (regs_regs_2_lpi_2[31:30])
      , (regs_regs_2_lpi_2[33:32]) , (regs_regs_2_lpi_2[35:34]) , (regs_regs_2_lpi_2[37:36])
      , (regs_regs_2_lpi_2[39:38]) , (regs_regs_2_lpi_2[41:40]) , (regs_regs_2_lpi_2[43:42])
      , (regs_regs_2_lpi_2[45:44]) , (regs_regs_2_lpi_2[47:46]) , (regs_regs_2_lpi_2[49:48])
      , (regs_regs_2_lpi_2[51:50]) , (regs_regs_2_lpi_2[53:52]) , (regs_regs_2_lpi_2[55:54])
      , (regs_regs_2_lpi_2[57:56]) , (regs_regs_2_lpi_2[59:58]) , (regs_regs_2_lpi_2[61:60])
      , (regs_regs_2_lpi_2[63:62]) , (regs_regs_2_lpi_2[65:64]) , (regs_regs_2_lpi_2[67:66])
      , (regs_regs_2_lpi_2[69:68]) , (regs_regs_2_lpi_2[71:70]) , (regs_regs_2_lpi_2[73:72])
      , (regs_regs_2_lpi_2[75:74]) , (regs_regs_2_lpi_2[77:76]) , (regs_regs_2_lpi_2[79:78])
      , (regs_regs_2_lpi_2[81:80]) , (regs_regs_2_lpi_2[83:82]) , (regs_regs_2_lpi_2[85:84])
      , (regs_regs_2_lpi_2[87:86]) , (regs_regs_2_lpi_2[89:88]) , (regs_regs_2_lpi_2[91:90])
      , (regs_regs_2_lpi_2[93:92]) , (regs_regs_2_lpi_2[95:94]) , (regs_regs_2_lpi_2[97:96])
      , (regs_regs_2_lpi_2[99:98]) , (regs_regs_2_lpi_2[101:100]) , (regs_regs_2_lpi_2[103:102])
      , (regs_regs_2_lpi_2[105:104]) , (regs_regs_2_lpi_2[107:106]) , (regs_regs_2_lpi_2[109:108])
      , (regs_regs_2_lpi_2[111:110]) , (regs_regs_2_lpi_2[113:112]) , (regs_regs_2_lpi_2[115:114])
      , (regs_regs_2_lpi_2[117:116]) , (regs_regs_2_lpi_2[119:118]) , (regs_regs_2_lpi_2[121:120])
      , (regs_regs_2_lpi_2[123:122]) , (regs_regs_2_lpi_2[125:124]) , (regs_regs_2_lpi_2[127:126])
      , (regs_regs_2_lpi_2[129:128]) , (regs_regs_2_lpi_2[131:130]) , (regs_regs_2_lpi_2[133:132])
      , (regs_regs_2_lpi_2[135:134]) , (regs_regs_2_lpi_2[137:136]) , (regs_regs_2_lpi_2[139:138])
      , (regs_regs_2_lpi_2[141:140]) , (regs_regs_2_lpi_2[143:142]) , (regs_regs_2_lpi_2[145:144])
      , (regs_regs_2_lpi_2[147:146]) , (regs_regs_2_lpi_2[149:148]) , (regs_regs_3_lpi_2[1:0])
      , (regs_regs_3_lpi_2[3:2]) , (regs_regs_3_lpi_2[5:4]) , (regs_regs_3_lpi_2[7:6])
      , (regs_regs_3_lpi_2[9:8]) , (regs_regs_3_lpi_2[11:10]) , (regs_regs_3_lpi_2[13:12])
      , (regs_regs_3_lpi_2[15:14]) , (regs_regs_3_lpi_2[17:16]) , (regs_regs_3_lpi_2[19:18])
      , (regs_regs_3_lpi_2[21:20]) , (regs_regs_3_lpi_2[23:22]) , (regs_regs_3_lpi_2[25:24])
      , (regs_regs_3_lpi_2[27:26]) , (regs_regs_3_lpi_2[29:28]) , (regs_regs_3_lpi_2[31:30])
      , (regs_regs_3_lpi_2[33:32]) , (regs_regs_3_lpi_2[35:34]) , (regs_regs_3_lpi_2[37:36])
      , (regs_regs_3_lpi_2[39:38]) , (regs_regs_3_lpi_2[41:40]) , (regs_regs_3_lpi_2[43:42])
      , (regs_regs_3_lpi_2[45:44]) , (regs_regs_3_lpi_2[47:46]) , (regs_regs_3_lpi_2[49:48])
      , (regs_regs_3_lpi_2[51:50]) , (regs_regs_3_lpi_2[53:52]) , (regs_regs_3_lpi_2[55:54])
      , (regs_regs_3_lpi_2[57:56]) , (regs_regs_3_lpi_2[59:58]) , (regs_regs_3_lpi_2[61:60])
      , (regs_regs_3_lpi_2[63:62]) , (regs_regs_3_lpi_2[65:64]) , (regs_regs_3_lpi_2[67:66])
      , (regs_regs_3_lpi_2[69:68]) , (regs_regs_3_lpi_2[71:70]) , (regs_regs_3_lpi_2[73:72])
      , (regs_regs_3_lpi_2[75:74]) , (regs_regs_3_lpi_2[77:76]) , (regs_regs_3_lpi_2[79:78])
      , (regs_regs_3_lpi_2[81:80]) , (regs_regs_3_lpi_2[83:82]) , (regs_regs_3_lpi_2[85:84])
      , (regs_regs_3_lpi_2[87:86]) , (regs_regs_3_lpi_2[89:88]) , (regs_regs_3_lpi_2[91:90])
      , (regs_regs_3_lpi_2[93:92]) , (regs_regs_3_lpi_2[95:94]) , (regs_regs_3_lpi_2[97:96])
      , (regs_regs_3_lpi_2[99:98]) , (regs_regs_3_lpi_2[101:100]) , (regs_regs_3_lpi_2[103:102])
      , (regs_regs_3_lpi_2[105:104]) , (regs_regs_3_lpi_2[107:106]) , (regs_regs_3_lpi_2[109:108])
      , (regs_regs_3_lpi_2[111:110]) , (regs_regs_3_lpi_2[113:112]) , (regs_regs_3_lpi_2[115:114])
      , (regs_regs_3_lpi_2[117:116]) , (regs_regs_3_lpi_2[119:118]) , (regs_regs_3_lpi_2[121:120])
      , (regs_regs_3_lpi_2[123:122]) , (regs_regs_3_lpi_2[125:124]) , (regs_regs_3_lpi_2[127:126])
      , (regs_regs_3_lpi_2[129:128]) , (regs_regs_3_lpi_2[131:130]) , (regs_regs_3_lpi_2[133:132])
      , (regs_regs_3_lpi_2[135:134]) , (regs_regs_3_lpi_2[137:136]) , (regs_regs_3_lpi_2[139:138])
      , (regs_regs_3_lpi_2[141:140]) , (regs_regs_3_lpi_2[143:142]) , (regs_regs_3_lpi_2[145:144])
      , (regs_regs_3_lpi_2[147:146]) , (regs_regs_3_lpi_2[149:148]) , (regs_regs_4_lpi_2[1:0])
      , (regs_regs_4_lpi_2[3:2]) , (regs_regs_4_lpi_2[5:4]) , (regs_regs_4_lpi_2[7:6])
      , (regs_regs_4_lpi_2[9:8]) , (regs_regs_4_lpi_2[11:10]) , (regs_regs_4_lpi_2[13:12])
      , (regs_regs_4_lpi_2[15:14]) , (regs_regs_4_lpi_2[17:16]) , (regs_regs_4_lpi_2[19:18])
      , (regs_regs_4_lpi_2[21:20]) , (regs_regs_4_lpi_2[23:22]) , (regs_regs_4_lpi_2[25:24])
      , (regs_regs_4_lpi_2[27:26]) , (regs_regs_4_lpi_2[29:28]) , (regs_regs_4_lpi_2[31:30])
      , (regs_regs_4_lpi_2[33:32]) , (regs_regs_4_lpi_2[35:34]) , (regs_regs_4_lpi_2[37:36])
      , (regs_regs_4_lpi_2[39:38]) , (regs_regs_4_lpi_2[41:40]) , (regs_regs_4_lpi_2[43:42])
      , (regs_regs_4_lpi_2[45:44]) , (regs_regs_4_lpi_2[47:46]) , (regs_regs_4_lpi_2[49:48])
      , (regs_regs_4_lpi_2[51:50]) , (regs_regs_4_lpi_2[53:52]) , (regs_regs_4_lpi_2[55:54])
      , (regs_regs_4_lpi_2[57:56]) , (regs_regs_4_lpi_2[59:58]) , (regs_regs_4_lpi_2[61:60])
      , (regs_regs_4_lpi_2[63:62]) , (regs_regs_4_lpi_2[65:64]) , (regs_regs_4_lpi_2[67:66])
      , (regs_regs_4_lpi_2[69:68]) , (regs_regs_4_lpi_2[71:70]) , (regs_regs_4_lpi_2[73:72])
      , (regs_regs_4_lpi_2[75:74]) , (regs_regs_4_lpi_2[77:76]) , (regs_regs_4_lpi_2[79:78])
      , (regs_regs_4_lpi_2[81:80]) , (regs_regs_4_lpi_2[83:82]) , (regs_regs_4_lpi_2[85:84])
      , (regs_regs_4_lpi_2[87:86]) , (regs_regs_4_lpi_2[89:88]) , (regs_regs_4_lpi_2[91:90])
      , (regs_regs_4_lpi_2[93:92]) , (regs_regs_4_lpi_2[95:94]) , (regs_regs_4_lpi_2[97:96])
      , (regs_regs_4_lpi_2[99:98]) , (regs_regs_4_lpi_2[101:100]) , (regs_regs_4_lpi_2[103:102])
      , (regs_regs_4_lpi_2[105:104]) , (regs_regs_4_lpi_2[107:106]) , (regs_regs_4_lpi_2[109:108])
      , (regs_regs_4_lpi_2[111:110]) , (regs_regs_4_lpi_2[113:112]) , (regs_regs_4_lpi_2[115:114])
      , (regs_regs_4_lpi_2[117:116]) , (regs_regs_4_lpi_2[119:118]) , (regs_regs_4_lpi_2[121:120])
      , (regs_regs_4_lpi_2[123:122]) , (regs_regs_4_lpi_2[125:124]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_sg1 = MUX_v_2_512_2({(regs_regs_0_lpi_2[3:2]) , (regs_regs_0_lpi_2[5:4])
      , (regs_regs_0_lpi_2[7:6]) , (regs_regs_0_lpi_2[9:8]) , (regs_regs_0_lpi_2[11:10])
      , (regs_regs_0_lpi_2[13:12]) , (regs_regs_0_lpi_2[15:14]) , (regs_regs_0_lpi_2[17:16])
      , (regs_regs_0_lpi_2[19:18]) , (regs_regs_0_lpi_2[21:20]) , (regs_regs_0_lpi_2[23:22])
      , (regs_regs_0_lpi_2[25:24]) , (regs_regs_0_lpi_2[27:26]) , (regs_regs_0_lpi_2[29:28])
      , (regs_regs_0_lpi_2[31:30]) , (regs_regs_0_lpi_2[33:32]) , (regs_regs_0_lpi_2[35:34])
      , (regs_regs_0_lpi_2[37:36]) , (regs_regs_0_lpi_2[39:38]) , (regs_regs_0_lpi_2[41:40])
      , (regs_regs_0_lpi_2[43:42]) , (regs_regs_0_lpi_2[45:44]) , (regs_regs_0_lpi_2[47:46])
      , (regs_regs_0_lpi_2[49:48]) , (regs_regs_0_lpi_2[51:50]) , (regs_regs_0_lpi_2[53:52])
      , (regs_regs_0_lpi_2[55:54]) , (regs_regs_0_lpi_2[57:56]) , (regs_regs_0_lpi_2[59:58])
      , (regs_regs_0_lpi_2[61:60]) , (regs_regs_0_lpi_2[63:62]) , (regs_regs_0_lpi_2[65:64])
      , (regs_regs_0_lpi_2[67:66]) , (regs_regs_0_lpi_2[69:68]) , (regs_regs_0_lpi_2[71:70])
      , (regs_regs_0_lpi_2[73:72]) , (regs_regs_0_lpi_2[75:74]) , (regs_regs_0_lpi_2[77:76])
      , (regs_regs_0_lpi_2[79:78]) , (regs_regs_0_lpi_2[81:80]) , (regs_regs_0_lpi_2[83:82])
      , (regs_regs_0_lpi_2[85:84]) , (regs_regs_0_lpi_2[87:86]) , (regs_regs_0_lpi_2[89:88])
      , (regs_regs_0_lpi_2[91:90]) , (regs_regs_0_lpi_2[93:92]) , (regs_regs_0_lpi_2[95:94])
      , (regs_regs_0_lpi_2[97:96]) , (regs_regs_0_lpi_2[99:98]) , (regs_regs_0_lpi_2[101:100])
      , (regs_regs_0_lpi_2[103:102]) , (regs_regs_0_lpi_2[105:104]) , (regs_regs_0_lpi_2[107:106])
      , (regs_regs_0_lpi_2[109:108]) , (regs_regs_0_lpi_2[111:110]) , (regs_regs_0_lpi_2[113:112])
      , (regs_regs_0_lpi_2[115:114]) , (regs_regs_0_lpi_2[117:116]) , (regs_regs_0_lpi_2[119:118])
      , (regs_regs_0_lpi_2[121:120]) , (regs_regs_0_lpi_2[123:122]) , (regs_regs_0_lpi_2[125:124])
      , (regs_regs_0_lpi_2[127:126]) , (regs_regs_0_lpi_2[129:128]) , (regs_regs_0_lpi_2[131:130])
      , (regs_regs_0_lpi_2[133:132]) , (regs_regs_0_lpi_2[135:134]) , (regs_regs_0_lpi_2[137:136])
      , (regs_regs_0_lpi_2[139:138]) , (regs_regs_0_lpi_2[141:140]) , (regs_regs_0_lpi_2[143:142])
      , (regs_regs_0_lpi_2[145:144]) , (regs_regs_0_lpi_2[147:146]) , (regs_regs_0_lpi_2[149:148])
      , (regs_regs_1_lpi_2[1:0]) , (regs_regs_1_lpi_2[3:2]) , (regs_regs_1_lpi_2[5:4])
      , (regs_regs_1_lpi_2[7:6]) , (regs_regs_1_lpi_2[9:8]) , (regs_regs_1_lpi_2[11:10])
      , (regs_regs_1_lpi_2[13:12]) , (regs_regs_1_lpi_2[15:14]) , (regs_regs_1_lpi_2[17:16])
      , (regs_regs_1_lpi_2[19:18]) , (regs_regs_1_lpi_2[21:20]) , (regs_regs_1_lpi_2[23:22])
      , (regs_regs_1_lpi_2[25:24]) , (regs_regs_1_lpi_2[27:26]) , (regs_regs_1_lpi_2[29:28])
      , (regs_regs_1_lpi_2[31:30]) , (regs_regs_1_lpi_2[33:32]) , (regs_regs_1_lpi_2[35:34])
      , (regs_regs_1_lpi_2[37:36]) , (regs_regs_1_lpi_2[39:38]) , (regs_regs_1_lpi_2[41:40])
      , (regs_regs_1_lpi_2[43:42]) , (regs_regs_1_lpi_2[45:44]) , (regs_regs_1_lpi_2[47:46])
      , (regs_regs_1_lpi_2[49:48]) , (regs_regs_1_lpi_2[51:50]) , (regs_regs_1_lpi_2[53:52])
      , (regs_regs_1_lpi_2[55:54]) , (regs_regs_1_lpi_2[57:56]) , (regs_regs_1_lpi_2[59:58])
      , (regs_regs_1_lpi_2[61:60]) , (regs_regs_1_lpi_2[63:62]) , (regs_regs_1_lpi_2[65:64])
      , (regs_regs_1_lpi_2[67:66]) , (regs_regs_1_lpi_2[69:68]) , (regs_regs_1_lpi_2[71:70])
      , (regs_regs_1_lpi_2[73:72]) , (regs_regs_1_lpi_2[75:74]) , (regs_regs_1_lpi_2[77:76])
      , (regs_regs_1_lpi_2[79:78]) , (regs_regs_1_lpi_2[81:80]) , (regs_regs_1_lpi_2[83:82])
      , (regs_regs_1_lpi_2[85:84]) , (regs_regs_1_lpi_2[87:86]) , (regs_regs_1_lpi_2[89:88])
      , (regs_regs_1_lpi_2[91:90]) , (regs_regs_1_lpi_2[93:92]) , (regs_regs_1_lpi_2[95:94])
      , (regs_regs_1_lpi_2[97:96]) , (regs_regs_1_lpi_2[99:98]) , (regs_regs_1_lpi_2[101:100])
      , (regs_regs_1_lpi_2[103:102]) , (regs_regs_1_lpi_2[105:104]) , (regs_regs_1_lpi_2[107:106])
      , (regs_regs_1_lpi_2[109:108]) , (regs_regs_1_lpi_2[111:110]) , (regs_regs_1_lpi_2[113:112])
      , (regs_regs_1_lpi_2[115:114]) , (regs_regs_1_lpi_2[117:116]) , (regs_regs_1_lpi_2[119:118])
      , (regs_regs_1_lpi_2[121:120]) , (regs_regs_1_lpi_2[123:122]) , (regs_regs_1_lpi_2[125:124])
      , (regs_regs_1_lpi_2[127:126]) , (regs_regs_1_lpi_2[129:128]) , (regs_regs_1_lpi_2[131:130])
      , (regs_regs_1_lpi_2[133:132]) , (regs_regs_1_lpi_2[135:134]) , (regs_regs_1_lpi_2[137:136])
      , (regs_regs_1_lpi_2[139:138]) , (regs_regs_1_lpi_2[141:140]) , (regs_regs_1_lpi_2[143:142])
      , (regs_regs_1_lpi_2[145:144]) , (regs_regs_1_lpi_2[147:146]) , (regs_regs_1_lpi_2[149:148])
      , (regs_regs_2_lpi_2[1:0]) , (regs_regs_2_lpi_2[3:2]) , (regs_regs_2_lpi_2[5:4])
      , (regs_regs_2_lpi_2[7:6]) , (regs_regs_2_lpi_2[9:8]) , (regs_regs_2_lpi_2[11:10])
      , (regs_regs_2_lpi_2[13:12]) , (regs_regs_2_lpi_2[15:14]) , (regs_regs_2_lpi_2[17:16])
      , (regs_regs_2_lpi_2[19:18]) , (regs_regs_2_lpi_2[21:20]) , (regs_regs_2_lpi_2[23:22])
      , (regs_regs_2_lpi_2[25:24]) , (regs_regs_2_lpi_2[27:26]) , (regs_regs_2_lpi_2[29:28])
      , (regs_regs_2_lpi_2[31:30]) , (regs_regs_2_lpi_2[33:32]) , (regs_regs_2_lpi_2[35:34])
      , (regs_regs_2_lpi_2[37:36]) , (regs_regs_2_lpi_2[39:38]) , (regs_regs_2_lpi_2[41:40])
      , (regs_regs_2_lpi_2[43:42]) , (regs_regs_2_lpi_2[45:44]) , (regs_regs_2_lpi_2[47:46])
      , (regs_regs_2_lpi_2[49:48]) , (regs_regs_2_lpi_2[51:50]) , (regs_regs_2_lpi_2[53:52])
      , (regs_regs_2_lpi_2[55:54]) , (regs_regs_2_lpi_2[57:56]) , (regs_regs_2_lpi_2[59:58])
      , (regs_regs_2_lpi_2[61:60]) , (regs_regs_2_lpi_2[63:62]) , (regs_regs_2_lpi_2[65:64])
      , (regs_regs_2_lpi_2[67:66]) , (regs_regs_2_lpi_2[69:68]) , (regs_regs_2_lpi_2[71:70])
      , (regs_regs_2_lpi_2[73:72]) , (regs_regs_2_lpi_2[75:74]) , (regs_regs_2_lpi_2[77:76])
      , (regs_regs_2_lpi_2[79:78]) , (regs_regs_2_lpi_2[81:80]) , (regs_regs_2_lpi_2[83:82])
      , (regs_regs_2_lpi_2[85:84]) , (regs_regs_2_lpi_2[87:86]) , (regs_regs_2_lpi_2[89:88])
      , (regs_regs_2_lpi_2[91:90]) , (regs_regs_2_lpi_2[93:92]) , (regs_regs_2_lpi_2[95:94])
      , (regs_regs_2_lpi_2[97:96]) , (regs_regs_2_lpi_2[99:98]) , (regs_regs_2_lpi_2[101:100])
      , (regs_regs_2_lpi_2[103:102]) , (regs_regs_2_lpi_2[105:104]) , (regs_regs_2_lpi_2[107:106])
      , (regs_regs_2_lpi_2[109:108]) , (regs_regs_2_lpi_2[111:110]) , (regs_regs_2_lpi_2[113:112])
      , (regs_regs_2_lpi_2[115:114]) , (regs_regs_2_lpi_2[117:116]) , (regs_regs_2_lpi_2[119:118])
      , (regs_regs_2_lpi_2[121:120]) , (regs_regs_2_lpi_2[123:122]) , (regs_regs_2_lpi_2[125:124])
      , (regs_regs_2_lpi_2[127:126]) , (regs_regs_2_lpi_2[129:128]) , (regs_regs_2_lpi_2[131:130])
      , (regs_regs_2_lpi_2[133:132]) , (regs_regs_2_lpi_2[135:134]) , (regs_regs_2_lpi_2[137:136])
      , (regs_regs_2_lpi_2[139:138]) , (regs_regs_2_lpi_2[141:140]) , (regs_regs_2_lpi_2[143:142])
      , (regs_regs_2_lpi_2[145:144]) , (regs_regs_2_lpi_2[147:146]) , (regs_regs_2_lpi_2[149:148])
      , (regs_regs_3_lpi_2[1:0]) , (regs_regs_3_lpi_2[3:2]) , (regs_regs_3_lpi_2[5:4])
      , (regs_regs_3_lpi_2[7:6]) , (regs_regs_3_lpi_2[9:8]) , (regs_regs_3_lpi_2[11:10])
      , (regs_regs_3_lpi_2[13:12]) , (regs_regs_3_lpi_2[15:14]) , (regs_regs_3_lpi_2[17:16])
      , (regs_regs_3_lpi_2[19:18]) , (regs_regs_3_lpi_2[21:20]) , (regs_regs_3_lpi_2[23:22])
      , (regs_regs_3_lpi_2[25:24]) , (regs_regs_3_lpi_2[27:26]) , (regs_regs_3_lpi_2[29:28])
      , (regs_regs_3_lpi_2[31:30]) , (regs_regs_3_lpi_2[33:32]) , (regs_regs_3_lpi_2[35:34])
      , (regs_regs_3_lpi_2[37:36]) , (regs_regs_3_lpi_2[39:38]) , (regs_regs_3_lpi_2[41:40])
      , (regs_regs_3_lpi_2[43:42]) , (regs_regs_3_lpi_2[45:44]) , (regs_regs_3_lpi_2[47:46])
      , (regs_regs_3_lpi_2[49:48]) , (regs_regs_3_lpi_2[51:50]) , (regs_regs_3_lpi_2[53:52])
      , (regs_regs_3_lpi_2[55:54]) , (regs_regs_3_lpi_2[57:56]) , (regs_regs_3_lpi_2[59:58])
      , (regs_regs_3_lpi_2[61:60]) , (regs_regs_3_lpi_2[63:62]) , (regs_regs_3_lpi_2[65:64])
      , (regs_regs_3_lpi_2[67:66]) , (regs_regs_3_lpi_2[69:68]) , (regs_regs_3_lpi_2[71:70])
      , (regs_regs_3_lpi_2[73:72]) , (regs_regs_3_lpi_2[75:74]) , (regs_regs_3_lpi_2[77:76])
      , (regs_regs_3_lpi_2[79:78]) , (regs_regs_3_lpi_2[81:80]) , (regs_regs_3_lpi_2[83:82])
      , (regs_regs_3_lpi_2[85:84]) , (regs_regs_3_lpi_2[87:86]) , (regs_regs_3_lpi_2[89:88])
      , (regs_regs_3_lpi_2[91:90]) , (regs_regs_3_lpi_2[93:92]) , (regs_regs_3_lpi_2[95:94])
      , (regs_regs_3_lpi_2[97:96]) , (regs_regs_3_lpi_2[99:98]) , (regs_regs_3_lpi_2[101:100])
      , (regs_regs_3_lpi_2[103:102]) , (regs_regs_3_lpi_2[105:104]) , (regs_regs_3_lpi_2[107:106])
      , (regs_regs_3_lpi_2[109:108]) , (regs_regs_3_lpi_2[111:110]) , (regs_regs_3_lpi_2[113:112])
      , (regs_regs_3_lpi_2[115:114]) , (regs_regs_3_lpi_2[117:116]) , (regs_regs_3_lpi_2[119:118])
      , (regs_regs_3_lpi_2[121:120]) , (regs_regs_3_lpi_2[123:122]) , (regs_regs_3_lpi_2[125:124])
      , (regs_regs_3_lpi_2[127:126]) , (regs_regs_3_lpi_2[129:128]) , (regs_regs_3_lpi_2[131:130])
      , (regs_regs_3_lpi_2[133:132]) , (regs_regs_3_lpi_2[135:134]) , (regs_regs_3_lpi_2[137:136])
      , (regs_regs_3_lpi_2[139:138]) , (regs_regs_3_lpi_2[141:140]) , (regs_regs_3_lpi_2[143:142])
      , (regs_regs_3_lpi_2[145:144]) , (regs_regs_3_lpi_2[147:146]) , (regs_regs_3_lpi_2[149:148])
      , (regs_regs_4_lpi_2[1:0]) , (regs_regs_4_lpi_2[3:2]) , (regs_regs_4_lpi_2[5:4])
      , (regs_regs_4_lpi_2[7:6]) , (regs_regs_4_lpi_2[9:8]) , (regs_regs_4_lpi_2[11:10])
      , (regs_regs_4_lpi_2[13:12]) , (regs_regs_4_lpi_2[15:14]) , (regs_regs_4_lpi_2[17:16])
      , (regs_regs_4_lpi_2[19:18]) , (regs_regs_4_lpi_2[21:20]) , (regs_regs_4_lpi_2[23:22])
      , (regs_regs_4_lpi_2[25:24]) , (regs_regs_4_lpi_2[27:26]) , (regs_regs_4_lpi_2[29:28])
      , (regs_regs_4_lpi_2[31:30]) , (regs_regs_4_lpi_2[33:32]) , (regs_regs_4_lpi_2[35:34])
      , (regs_regs_4_lpi_2[37:36]) , (regs_regs_4_lpi_2[39:38]) , (regs_regs_4_lpi_2[41:40])
      , (regs_regs_4_lpi_2[43:42]) , (regs_regs_4_lpi_2[45:44]) , (regs_regs_4_lpi_2[47:46])
      , (regs_regs_4_lpi_2[49:48]) , (regs_regs_4_lpi_2[51:50]) , (regs_regs_4_lpi_2[53:52])
      , (regs_regs_4_lpi_2[55:54]) , (regs_regs_4_lpi_2[57:56]) , (regs_regs_4_lpi_2[59:58])
      , (regs_regs_4_lpi_2[61:60]) , (regs_regs_4_lpi_2[63:62]) , (regs_regs_4_lpi_2[65:64])
      , (regs_regs_4_lpi_2[67:66]) , (regs_regs_4_lpi_2[69:68]) , (regs_regs_4_lpi_2[71:70])
      , (regs_regs_4_lpi_2[73:72]) , (regs_regs_4_lpi_2[75:74]) , (regs_regs_4_lpi_2[77:76])
      , (regs_regs_4_lpi_2[79:78]) , (regs_regs_4_lpi_2[81:80]) , (regs_regs_4_lpi_2[83:82])
      , (regs_regs_4_lpi_2[85:84]) , (regs_regs_4_lpi_2[87:86]) , (regs_regs_4_lpi_2[89:88])
      , (regs_regs_4_lpi_2[91:90]) , (regs_regs_4_lpi_2[93:92]) , (regs_regs_4_lpi_2[95:94])
      , (regs_regs_4_lpi_2[97:96]) , (regs_regs_4_lpi_2[99:98]) , (regs_regs_4_lpi_2[101:100])
      , (regs_regs_4_lpi_2[103:102]) , (regs_regs_4_lpi_2[105:104]) , (regs_regs_4_lpi_2[107:106])
      , (regs_regs_4_lpi_2[109:108]) , (regs_regs_4_lpi_2[111:110]) , (regs_regs_4_lpi_2[113:112])
      , (regs_regs_4_lpi_2[115:114]) , (regs_regs_4_lpi_2[117:116]) , (regs_regs_4_lpi_2[119:118])
      , (regs_regs_4_lpi_2[121:120]) , (regs_regs_4_lpi_2[123:122]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign ACC1_for_slc_1_svs_1 = MUX_v_2_512_2({(regs_regs_0_lpi_2[1:0]) , (regs_regs_0_lpi_2[3:2])
      , (regs_regs_0_lpi_2[5:4]) , (regs_regs_0_lpi_2[7:6]) , (regs_regs_0_lpi_2[9:8])
      , (regs_regs_0_lpi_2[11:10]) , (regs_regs_0_lpi_2[13:12]) , (regs_regs_0_lpi_2[15:14])
      , (regs_regs_0_lpi_2[17:16]) , (regs_regs_0_lpi_2[19:18]) , (regs_regs_0_lpi_2[21:20])
      , (regs_regs_0_lpi_2[23:22]) , (regs_regs_0_lpi_2[25:24]) , (regs_regs_0_lpi_2[27:26])
      , (regs_regs_0_lpi_2[29:28]) , (regs_regs_0_lpi_2[31:30]) , (regs_regs_0_lpi_2[33:32])
      , (regs_regs_0_lpi_2[35:34]) , (regs_regs_0_lpi_2[37:36]) , (regs_regs_0_lpi_2[39:38])
      , (regs_regs_0_lpi_2[41:40]) , (regs_regs_0_lpi_2[43:42]) , (regs_regs_0_lpi_2[45:44])
      , (regs_regs_0_lpi_2[47:46]) , (regs_regs_0_lpi_2[49:48]) , (regs_regs_0_lpi_2[51:50])
      , (regs_regs_0_lpi_2[53:52]) , (regs_regs_0_lpi_2[55:54]) , (regs_regs_0_lpi_2[57:56])
      , (regs_regs_0_lpi_2[59:58]) , (regs_regs_0_lpi_2[61:60]) , (regs_regs_0_lpi_2[63:62])
      , (regs_regs_0_lpi_2[65:64]) , (regs_regs_0_lpi_2[67:66]) , (regs_regs_0_lpi_2[69:68])
      , (regs_regs_0_lpi_2[71:70]) , (regs_regs_0_lpi_2[73:72]) , (regs_regs_0_lpi_2[75:74])
      , (regs_regs_0_lpi_2[77:76]) , (regs_regs_0_lpi_2[79:78]) , (regs_regs_0_lpi_2[81:80])
      , (regs_regs_0_lpi_2[83:82]) , (regs_regs_0_lpi_2[85:84]) , (regs_regs_0_lpi_2[87:86])
      , (regs_regs_0_lpi_2[89:88]) , (regs_regs_0_lpi_2[91:90]) , (regs_regs_0_lpi_2[93:92])
      , (regs_regs_0_lpi_2[95:94]) , (regs_regs_0_lpi_2[97:96]) , (regs_regs_0_lpi_2[99:98])
      , (regs_regs_0_lpi_2[101:100]) , (regs_regs_0_lpi_2[103:102]) , (regs_regs_0_lpi_2[105:104])
      , (regs_regs_0_lpi_2[107:106]) , (regs_regs_0_lpi_2[109:108]) , (regs_regs_0_lpi_2[111:110])
      , (regs_regs_0_lpi_2[113:112]) , (regs_regs_0_lpi_2[115:114]) , (regs_regs_0_lpi_2[117:116])
      , (regs_regs_0_lpi_2[119:118]) , (regs_regs_0_lpi_2[121:120]) , (regs_regs_0_lpi_2[123:122])
      , (regs_regs_0_lpi_2[125:124]) , (regs_regs_0_lpi_2[127:126]) , (regs_regs_0_lpi_2[129:128])
      , (regs_regs_0_lpi_2[131:130]) , (regs_regs_0_lpi_2[133:132]) , (regs_regs_0_lpi_2[135:134])
      , (regs_regs_0_lpi_2[137:136]) , (regs_regs_0_lpi_2[139:138]) , (regs_regs_0_lpi_2[141:140])
      , (regs_regs_0_lpi_2[143:142]) , (regs_regs_0_lpi_2[145:144]) , (regs_regs_0_lpi_2[147:146])
      , (regs_regs_0_lpi_2[149:148]) , (regs_regs_1_lpi_2[1:0]) , (regs_regs_1_lpi_2[3:2])
      , (regs_regs_1_lpi_2[5:4]) , (regs_regs_1_lpi_2[7:6]) , (regs_regs_1_lpi_2[9:8])
      , (regs_regs_1_lpi_2[11:10]) , (regs_regs_1_lpi_2[13:12]) , (regs_regs_1_lpi_2[15:14])
      , (regs_regs_1_lpi_2[17:16]) , (regs_regs_1_lpi_2[19:18]) , (regs_regs_1_lpi_2[21:20])
      , (regs_regs_1_lpi_2[23:22]) , (regs_regs_1_lpi_2[25:24]) , (regs_regs_1_lpi_2[27:26])
      , (regs_regs_1_lpi_2[29:28]) , (regs_regs_1_lpi_2[31:30]) , (regs_regs_1_lpi_2[33:32])
      , (regs_regs_1_lpi_2[35:34]) , (regs_regs_1_lpi_2[37:36]) , (regs_regs_1_lpi_2[39:38])
      , (regs_regs_1_lpi_2[41:40]) , (regs_regs_1_lpi_2[43:42]) , (regs_regs_1_lpi_2[45:44])
      , (regs_regs_1_lpi_2[47:46]) , (regs_regs_1_lpi_2[49:48]) , (regs_regs_1_lpi_2[51:50])
      , (regs_regs_1_lpi_2[53:52]) , (regs_regs_1_lpi_2[55:54]) , (regs_regs_1_lpi_2[57:56])
      , (regs_regs_1_lpi_2[59:58]) , (regs_regs_1_lpi_2[61:60]) , (regs_regs_1_lpi_2[63:62])
      , (regs_regs_1_lpi_2[65:64]) , (regs_regs_1_lpi_2[67:66]) , (regs_regs_1_lpi_2[69:68])
      , (regs_regs_1_lpi_2[71:70]) , (regs_regs_1_lpi_2[73:72]) , (regs_regs_1_lpi_2[75:74])
      , (regs_regs_1_lpi_2[77:76]) , (regs_regs_1_lpi_2[79:78]) , (regs_regs_1_lpi_2[81:80])
      , (regs_regs_1_lpi_2[83:82]) , (regs_regs_1_lpi_2[85:84]) , (regs_regs_1_lpi_2[87:86])
      , (regs_regs_1_lpi_2[89:88]) , (regs_regs_1_lpi_2[91:90]) , (regs_regs_1_lpi_2[93:92])
      , (regs_regs_1_lpi_2[95:94]) , (regs_regs_1_lpi_2[97:96]) , (regs_regs_1_lpi_2[99:98])
      , (regs_regs_1_lpi_2[101:100]) , (regs_regs_1_lpi_2[103:102]) , (regs_regs_1_lpi_2[105:104])
      , (regs_regs_1_lpi_2[107:106]) , (regs_regs_1_lpi_2[109:108]) , (regs_regs_1_lpi_2[111:110])
      , (regs_regs_1_lpi_2[113:112]) , (regs_regs_1_lpi_2[115:114]) , (regs_regs_1_lpi_2[117:116])
      , (regs_regs_1_lpi_2[119:118]) , (regs_regs_1_lpi_2[121:120]) , (regs_regs_1_lpi_2[123:122])
      , (regs_regs_1_lpi_2[125:124]) , (regs_regs_1_lpi_2[127:126]) , (regs_regs_1_lpi_2[129:128])
      , (regs_regs_1_lpi_2[131:130]) , (regs_regs_1_lpi_2[133:132]) , (regs_regs_1_lpi_2[135:134])
      , (regs_regs_1_lpi_2[137:136]) , (regs_regs_1_lpi_2[139:138]) , (regs_regs_1_lpi_2[141:140])
      , (regs_regs_1_lpi_2[143:142]) , (regs_regs_1_lpi_2[145:144]) , (regs_regs_1_lpi_2[147:146])
      , (regs_regs_1_lpi_2[149:148]) , (regs_regs_2_lpi_2[1:0]) , (regs_regs_2_lpi_2[3:2])
      , (regs_regs_2_lpi_2[5:4]) , (regs_regs_2_lpi_2[7:6]) , (regs_regs_2_lpi_2[9:8])
      , (regs_regs_2_lpi_2[11:10]) , (regs_regs_2_lpi_2[13:12]) , (regs_regs_2_lpi_2[15:14])
      , (regs_regs_2_lpi_2[17:16]) , (regs_regs_2_lpi_2[19:18]) , (regs_regs_2_lpi_2[21:20])
      , (regs_regs_2_lpi_2[23:22]) , (regs_regs_2_lpi_2[25:24]) , (regs_regs_2_lpi_2[27:26])
      , (regs_regs_2_lpi_2[29:28]) , (regs_regs_2_lpi_2[31:30]) , (regs_regs_2_lpi_2[33:32])
      , (regs_regs_2_lpi_2[35:34]) , (regs_regs_2_lpi_2[37:36]) , (regs_regs_2_lpi_2[39:38])
      , (regs_regs_2_lpi_2[41:40]) , (regs_regs_2_lpi_2[43:42]) , (regs_regs_2_lpi_2[45:44])
      , (regs_regs_2_lpi_2[47:46]) , (regs_regs_2_lpi_2[49:48]) , (regs_regs_2_lpi_2[51:50])
      , (regs_regs_2_lpi_2[53:52]) , (regs_regs_2_lpi_2[55:54]) , (regs_regs_2_lpi_2[57:56])
      , (regs_regs_2_lpi_2[59:58]) , (regs_regs_2_lpi_2[61:60]) , (regs_regs_2_lpi_2[63:62])
      , (regs_regs_2_lpi_2[65:64]) , (regs_regs_2_lpi_2[67:66]) , (regs_regs_2_lpi_2[69:68])
      , (regs_regs_2_lpi_2[71:70]) , (regs_regs_2_lpi_2[73:72]) , (regs_regs_2_lpi_2[75:74])
      , (regs_regs_2_lpi_2[77:76]) , (regs_regs_2_lpi_2[79:78]) , (regs_regs_2_lpi_2[81:80])
      , (regs_regs_2_lpi_2[83:82]) , (regs_regs_2_lpi_2[85:84]) , (regs_regs_2_lpi_2[87:86])
      , (regs_regs_2_lpi_2[89:88]) , (regs_regs_2_lpi_2[91:90]) , (regs_regs_2_lpi_2[93:92])
      , (regs_regs_2_lpi_2[95:94]) , (regs_regs_2_lpi_2[97:96]) , (regs_regs_2_lpi_2[99:98])
      , (regs_regs_2_lpi_2[101:100]) , (regs_regs_2_lpi_2[103:102]) , (regs_regs_2_lpi_2[105:104])
      , (regs_regs_2_lpi_2[107:106]) , (regs_regs_2_lpi_2[109:108]) , (regs_regs_2_lpi_2[111:110])
      , (regs_regs_2_lpi_2[113:112]) , (regs_regs_2_lpi_2[115:114]) , (regs_regs_2_lpi_2[117:116])
      , (regs_regs_2_lpi_2[119:118]) , (regs_regs_2_lpi_2[121:120]) , (regs_regs_2_lpi_2[123:122])
      , (regs_regs_2_lpi_2[125:124]) , (regs_regs_2_lpi_2[127:126]) , (regs_regs_2_lpi_2[129:128])
      , (regs_regs_2_lpi_2[131:130]) , (regs_regs_2_lpi_2[133:132]) , (regs_regs_2_lpi_2[135:134])
      , (regs_regs_2_lpi_2[137:136]) , (regs_regs_2_lpi_2[139:138]) , (regs_regs_2_lpi_2[141:140])
      , (regs_regs_2_lpi_2[143:142]) , (regs_regs_2_lpi_2[145:144]) , (regs_regs_2_lpi_2[147:146])
      , (regs_regs_2_lpi_2[149:148]) , (regs_regs_3_lpi_2[1:0]) , (regs_regs_3_lpi_2[3:2])
      , (regs_regs_3_lpi_2[5:4]) , (regs_regs_3_lpi_2[7:6]) , (regs_regs_3_lpi_2[9:8])
      , (regs_regs_3_lpi_2[11:10]) , (regs_regs_3_lpi_2[13:12]) , (regs_regs_3_lpi_2[15:14])
      , (regs_regs_3_lpi_2[17:16]) , (regs_regs_3_lpi_2[19:18]) , (regs_regs_3_lpi_2[21:20])
      , (regs_regs_3_lpi_2[23:22]) , (regs_regs_3_lpi_2[25:24]) , (regs_regs_3_lpi_2[27:26])
      , (regs_regs_3_lpi_2[29:28]) , (regs_regs_3_lpi_2[31:30]) , (regs_regs_3_lpi_2[33:32])
      , (regs_regs_3_lpi_2[35:34]) , (regs_regs_3_lpi_2[37:36]) , (regs_regs_3_lpi_2[39:38])
      , (regs_regs_3_lpi_2[41:40]) , (regs_regs_3_lpi_2[43:42]) , (regs_regs_3_lpi_2[45:44])
      , (regs_regs_3_lpi_2[47:46]) , (regs_regs_3_lpi_2[49:48]) , (regs_regs_3_lpi_2[51:50])
      , (regs_regs_3_lpi_2[53:52]) , (regs_regs_3_lpi_2[55:54]) , (regs_regs_3_lpi_2[57:56])
      , (regs_regs_3_lpi_2[59:58]) , (regs_regs_3_lpi_2[61:60]) , (regs_regs_3_lpi_2[63:62])
      , (regs_regs_3_lpi_2[65:64]) , (regs_regs_3_lpi_2[67:66]) , (regs_regs_3_lpi_2[69:68])
      , (regs_regs_3_lpi_2[71:70]) , (regs_regs_3_lpi_2[73:72]) , (regs_regs_3_lpi_2[75:74])
      , (regs_regs_3_lpi_2[77:76]) , (regs_regs_3_lpi_2[79:78]) , (regs_regs_3_lpi_2[81:80])
      , (regs_regs_3_lpi_2[83:82]) , (regs_regs_3_lpi_2[85:84]) , (regs_regs_3_lpi_2[87:86])
      , (regs_regs_3_lpi_2[89:88]) , (regs_regs_3_lpi_2[91:90]) , (regs_regs_3_lpi_2[93:92])
      , (regs_regs_3_lpi_2[95:94]) , (regs_regs_3_lpi_2[97:96]) , (regs_regs_3_lpi_2[99:98])
      , (regs_regs_3_lpi_2[101:100]) , (regs_regs_3_lpi_2[103:102]) , (regs_regs_3_lpi_2[105:104])
      , (regs_regs_3_lpi_2[107:106]) , (regs_regs_3_lpi_2[109:108]) , (regs_regs_3_lpi_2[111:110])
      , (regs_regs_3_lpi_2[113:112]) , (regs_regs_3_lpi_2[115:114]) , (regs_regs_3_lpi_2[117:116])
      , (regs_regs_3_lpi_2[119:118]) , (regs_regs_3_lpi_2[121:120]) , (regs_regs_3_lpi_2[123:122])
      , (regs_regs_3_lpi_2[125:124]) , (regs_regs_3_lpi_2[127:126]) , (regs_regs_3_lpi_2[129:128])
      , (regs_regs_3_lpi_2[131:130]) , (regs_regs_3_lpi_2[133:132]) , (regs_regs_3_lpi_2[135:134])
      , (regs_regs_3_lpi_2[137:136]) , (regs_regs_3_lpi_2[139:138]) , (regs_regs_3_lpi_2[141:140])
      , (regs_regs_3_lpi_2[143:142]) , (regs_regs_3_lpi_2[145:144]) , (regs_regs_3_lpi_2[147:146])
      , (regs_regs_3_lpi_2[149:148]) , (regs_regs_4_lpi_2[1:0]) , (regs_regs_4_lpi_2[3:2])
      , (regs_regs_4_lpi_2[5:4]) , (regs_regs_4_lpi_2[7:6]) , (regs_regs_4_lpi_2[9:8])
      , (regs_regs_4_lpi_2[11:10]) , (regs_regs_4_lpi_2[13:12]) , (regs_regs_4_lpi_2[15:14])
      , (regs_regs_4_lpi_2[17:16]) , (regs_regs_4_lpi_2[19:18]) , (regs_regs_4_lpi_2[21:20])
      , (regs_regs_4_lpi_2[23:22]) , (regs_regs_4_lpi_2[25:24]) , (regs_regs_4_lpi_2[27:26])
      , (regs_regs_4_lpi_2[29:28]) , (regs_regs_4_lpi_2[31:30]) , (regs_regs_4_lpi_2[33:32])
      , (regs_regs_4_lpi_2[35:34]) , (regs_regs_4_lpi_2[37:36]) , (regs_regs_4_lpi_2[39:38])
      , (regs_regs_4_lpi_2[41:40]) , (regs_regs_4_lpi_2[43:42]) , (regs_regs_4_lpi_2[45:44])
      , (regs_regs_4_lpi_2[47:46]) , (regs_regs_4_lpi_2[49:48]) , (regs_regs_4_lpi_2[51:50])
      , (regs_regs_4_lpi_2[53:52]) , (regs_regs_4_lpi_2[55:54]) , (regs_regs_4_lpi_2[57:56])
      , (regs_regs_4_lpi_2[59:58]) , (regs_regs_4_lpi_2[61:60]) , (regs_regs_4_lpi_2[63:62])
      , (regs_regs_4_lpi_2[65:64]) , (regs_regs_4_lpi_2[67:66]) , (regs_regs_4_lpi_2[69:68])
      , (regs_regs_4_lpi_2[71:70]) , (regs_regs_4_lpi_2[73:72]) , (regs_regs_4_lpi_2[75:74])
      , (regs_regs_4_lpi_2[77:76]) , (regs_regs_4_lpi_2[79:78]) , (regs_regs_4_lpi_2[81:80])
      , (regs_regs_4_lpi_2[83:82]) , (regs_regs_4_lpi_2[85:84]) , (regs_regs_4_lpi_2[87:86])
      , (regs_regs_4_lpi_2[89:88]) , (regs_regs_4_lpi_2[91:90]) , (regs_regs_4_lpi_2[93:92])
      , (regs_regs_4_lpi_2[95:94]) , (regs_regs_4_lpi_2[97:96]) , (regs_regs_4_lpi_2[99:98])
      , (regs_regs_4_lpi_2[101:100]) , (regs_regs_4_lpi_2[103:102]) , (regs_regs_4_lpi_2[105:104])
      , (regs_regs_4_lpi_2[107:106]) , (regs_regs_4_lpi_2[109:108]) , (regs_regs_4_lpi_2[111:110])
      , (regs_regs_4_lpi_2[113:112]) , (regs_regs_4_lpi_2[115:114]) , (regs_regs_4_lpi_2[117:116])
      , (regs_regs_4_lpi_2[119:118]) , (regs_regs_4_lpi_2[121:120]) , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0
      , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0 , 2'b0}, ACC1_for_if_acc_ssc);
  assign nl_ACC1_for_if_acc_ssc = conv_u2u_6_9(conv_s2u_4_6({1'b1 , (~ ACC1_for_j_1_lpi_2)})
      + ({(ACC1_for_j_1_lpi_2[1:0]) , 4'b1})) + conv_u2u_18_9(conv_u2u_3_9(i_1_lpi_2)
      * 9'b1001011);
  assign ACC1_for_if_acc_ssc = nl_ACC1_for_if_acc_ssc[8:0];
  assign SHIFT_i_1_lpi_2_dfm_2_mx0 = MUX_v_3_2_2({SHIFT_i_1_lpi_5 , 3'b100}, exit_ACC1_1_sva);
  assign exit_SHIFT_lpi_2_dfm_2 = exit_SHIFT_lpi_2 & (~ exit_ACC1_1_sva);
  assign SHIFT_and_8_cse = exit_ACC1_for_lpi_2_dfm_1_mx2 & exit_SHIFT_lpi_2_dfm_2;
  assign SHIFT_and_cse = (~ exit_ACC1_for_lpi_2_dfm_1_mx2) & exit_SHIFT_lpi_2_dfm_2;
  assign SHIFT_if_else_else_else_slc_regs_regs_ctmp_sva = MUX_v_150_4_2({regs_regs_0_lpi_2
      , regs_regs_1_lpi_2 , regs_regs_2_lpi_2 , regs_regs_3_lpi_2}, (SHIFT_i_1_lpi_2_dfm_2_mx0[1:0])
      + 2'b11);
  assign nl_SHIFT_acc_1_psp = SHIFT_i_1_lpi_2_dfm_2_mx0 + 3'b111;
  assign SHIFT_acc_1_psp = nl_SHIFT_acc_1_psp[2:0];
  assign SHIFT_mux_2_tmp = MUX_v_3_2_2({SHIFT_i_1_lpi_5 , 3'b100}, exit_ACC1_1_sva);
  assign and_dcpl = (~ ACC1_for_nand_tmp) & (ACC1_for_acc_itm[2]);
  assign or_dcpl_80 = (~ exit_SHIFT_lpi_2) | exit_ACC1_1_sva;
  assign or_dcpl_83 = exit_ACC1_1_sva | (ACC1_acc_itm[2]);
  assign or_dcpl_85 = and_dcpl | (~ exit_SHIFT_lpi_2);
  assign and_88_cse = exit_SHIFT_lpi_2_dfm_2 & FRAME_stage_0;
  assign and_89_cse = or_dcpl_80 & FRAME_stage_0;
  assign and_dcpl_90 = ~((SHIFT_mux_2_tmp[0]) | (SHIFT_mux_2_tmp[1]));
  assign or_dcpl_93 = exit_SHIFT_lpi_2_dfm_2 | (SHIFT_mux_2_tmp[0]);
  assign nor_8_cse = ~(exit_SHIFT_lpi_2_dfm_2 | (SHIFT_acc_1_psp[2]));
  assign or_dcpl_113 = nor_8_cse | SHIFT_and_cse;
  assign and_dcpl_136 = (~ exit_SHIFT_lpi_2_dfm_2) & (SHIFT_acc_1_psp[2]);
  assign or_dcpl_115 = (SHIFT_and_8_cse & ACC1_for_nand_tmp & (~ (ACC1_acc_itm[2])))
      | nor_8_cse;
  assign or_dcpl_116 = and_dcpl_136 | (SHIFT_and_8_cse & (ACC1_acc_itm[2]));
  always @(posedge clk or negedge arst_n) begin
    if ( ~ arst_n ) begin
      vout_rsc_mgc_out_stdreg_d <= 30'b0;
      FRAME_stage_0 <= 1'b0;
      FRAME_p_1_sva <= 19'b0;
      i_1_lpi_2 <= 3'b0;
      exit_ACC1_lpi_2 <= 1'b0;
      ACC1_for_j_1_lpi_2 <= 3'b0;
      regs_regs_4_lpi_2 <= 150'b0;
      regs_regs_3_lpi_2 <= 150'b0;
      regs_regs_2_lpi_2 <= 150'b0;
      regs_regs_1_lpi_2 <= 150'b0;
      regs_regs_0_lpi_2 <= 150'b0;
      exit_SHIFT_lpi_2 <= 1'b0;
      exit_ACC1_1_sva <= 1'b0;
      SHIFT_i_1_lpi_5 <= 3'b0;
      apply_lpi_2 <= 1'b0;
      exit_ACC1_for_lpi_2_dfm_1 <= 1'b0;
      regs_operator_din_lpi_2 <= 150'b0;
      apply_lpi_2_dfm_2 <= 1'b0;
      exit_SHIFT_lpi_2_dfm_1 <= 1'b0;
      ACC1_for_j_1_lpi_2_dfm_4 <= 3'b0;
      i_1_lpi_2_dfm_2 <= 3'b0;
      exit_ACC1_lpi_2_dfm_3 <= 1'b0;
      regs_regs_4_lpi_2_dfm_1 <= 150'b0;
      regs_regs_3_lpi_2_dfm_1 <= 150'b0;
      regs_regs_2_lpi_2_dfm_1 <= 150'b0;
      regs_regs_1_lpi_2_dfm_1 <= 150'b0;
      regs_regs_0_lpi_2_dfm_1 <= 150'b0;
    end
    else begin
      if ( en ) begin
        vout_rsc_mgc_out_stdreg_d <= (vout_rsc_mgc_out_stdreg_d & (signext_30_1(~(exit_SHIFT_lpi_2
            & (~ (ACC1_acc_itm[2])) & (fsm_output[1]) & FRAME_stage_0 & (~((~((~((ACC1_for_acc_itm[2])
            | apply_lpi_2)) | ACC1_for_nand_tmp)) | exit_ACC1_1_sva)))))) | (signext_30_1(exit_SHIFT_lpi_2_dfm_2
            & (~(ACC1_for_nand_tmp | (ACC1_for_acc_itm[2]))) & (~ (ACC1_acc_itm[2]))
            & (fsm_output[1]) & FRAME_stage_0 & apply_lpi_2));
        FRAME_stage_0 <= ~((~(FRAME_stage_0 & (or_dcpl_85 | or_dcpl_83 | (readslicef_8_1_7((conv_u2s_7_8(FRAME_p_1_sva_1[18:12])
            + 8'b10110101)))))) & (fsm_output[1]));
        FRAME_p_1_sva <= (MUX_v_19_2_2({FRAME_p_1_sva_1 , FRAME_p_1_sva}, or_dcpl_85
            | or_dcpl_83)) & (signext_19_1(fsm_output[1]));
        i_1_lpi_2 <= MUX1HOT_v_3_3_2({i_1_lpi_2 , i_1_lpi_2_dfm_2 , i_1_lpi_2_dfm_2_mx1w0},
            {(~ (fsm_output[1])) , and_151_cse , and_152_cse});
        exit_ACC1_lpi_2 <= MUX_s_1_2_2({exit_ACC1_lpi_2 , (MUX1HOT_s_1_3_2({exit_ACC1_lpi_2_dfm_1_mx0
            , (exit_ACC1_lpi_2 & (~ (SHIFT_acc_1_psp[2]))) , exit_ACC1_lpi_2_dfm_3},
            {and_88_cse , and_89_cse , (~ FRAME_stage_0)}))}, fsm_output[1]);
        ACC1_for_j_1_lpi_2 <= MUX1HOT_v_3_3_2({ACC1_for_j_1_lpi_2 , ACC1_for_j_1_lpi_2_dfm_4
            , ACC1_for_j_1_lpi_2_dfm_4_mx1w0}, {(~ (fsm_output[1])) , and_151_cse
            , and_152_cse});
        regs_regs_4_lpi_2 <= MUX1HOT_v_150_3_2({regs_regs_4_lpi_2 , SHIFT_if_else_else_else_slc_regs_regs_ctmp_sva
            , regs_regs_4_lpi_2_dfm_1}, {(~((fsm_output[1]) & (~((or_dcpl_93 | (SHIFT_mux_2_tmp[1])
            | (~ (SHIFT_mux_2_tmp[2]))) & FRAME_stage_0)))) , (and_89_cse & and_dcpl_90
            & (SHIFT_mux_2_tmp[2]) & (fsm_output[1])) , and_151_cse});
        regs_regs_3_lpi_2 <= MUX1HOT_v_150_3_2({regs_regs_3_lpi_2 , SHIFT_if_else_else_else_slc_regs_regs_ctmp_sva
            , regs_regs_3_lpi_2_dfm_1}, {(~((fsm_output[1]) & (~((exit_SHIFT_lpi_2_dfm_2
            | (~((SHIFT_mux_2_tmp[0]) & (SHIFT_mux_2_tmp[1])))) & FRAME_stage_0))))
            , (and_89_cse & (SHIFT_mux_2_tmp[0]) & (SHIFT_mux_2_tmp[1]) & (fsm_output[1]))
            , and_151_cse});
        regs_regs_2_lpi_2 <= MUX1HOT_v_150_3_2({regs_regs_2_lpi_2 , SHIFT_if_else_else_else_slc_regs_regs_ctmp_sva
            , regs_regs_2_lpi_2_dfm_1}, {(~((fsm_output[1]) & (~((exit_SHIFT_lpi_2_dfm_2
            | (SHIFT_mux_2_tmp[0]) | (~ (SHIFT_mux_2_tmp[1]))) & FRAME_stage_0))))
            , (and_89_cse & (~ (SHIFT_mux_2_tmp[0])) & (SHIFT_mux_2_tmp[1]) & (fsm_output[1]))
            , and_151_cse});
        regs_regs_1_lpi_2 <= MUX1HOT_v_150_3_2({regs_regs_1_lpi_2 , SHIFT_if_else_else_else_slc_regs_regs_ctmp_sva
            , regs_regs_1_lpi_2_dfm_1}, {(~((fsm_output[1]) & (~((exit_SHIFT_lpi_2_dfm_2
            | (~ (SHIFT_mux_2_tmp[0])) | (SHIFT_mux_2_tmp[1])) & FRAME_stage_0))))
            , (and_89_cse & (SHIFT_mux_2_tmp[0]) & (~ (SHIFT_mux_2_tmp[1])) & (fsm_output[1]))
            , and_151_cse});
        regs_regs_0_lpi_2 <= MUX1HOT_v_150_3_2({regs_regs_0_lpi_2 , regs_operator_din_lpi_2_mx0
            , regs_regs_0_lpi_2_dfm_1}, {(~((fsm_output[1]) & (~((or_dcpl_93 | (SHIFT_mux_2_tmp[1])
            | (SHIFT_mux_2_tmp[2])) & FRAME_stage_0)))) , (and_89_cse & and_dcpl_90
            & (~ (SHIFT_mux_2_tmp[2])) & (fsm_output[1])) , and_151_cse});
        exit_SHIFT_lpi_2 <= MUX_s_1_2_2({exit_SHIFT_lpi_2 , (MUX1HOT_s_1_3_2({exit_SHIFT_lpi_2_dfm_2
            , (SHIFT_acc_1_psp[2]) , exit_SHIFT_lpi_2_dfm_1}, {and_88_cse , and_89_cse
            , (~ FRAME_stage_0)}))}, fsm_output[1]);
        exit_ACC1_1_sva <= ~((~(((~ (ACC1_for_acc_itm[2])) | ACC1_for_nand_tmp) &
            exit_ACC1_lpi_2_dfm_1_mx0 & exit_SHIFT_lpi_2_dfm_2)) & (fsm_output[1]));
        SHIFT_i_1_lpi_5 <= MUX_v_3_2_2({SHIFT_acc_1_psp , SHIFT_i_1_lpi_5}, exit_SHIFT_lpi_2_dfm_2);
        apply_lpi_2 <= MUX_s_1_2_2({apply_lpi_2 , (MUX1HOT_s_1_3_2({apply_lpi_2_dfm_1
            , apply_lpi_2_dfm , apply_lpi_2_dfm_2}, {and_88_cse , and_89_cse , (~
            FRAME_stage_0)}))}, fsm_output[1]);
        exit_ACC1_for_lpi_2_dfm_1 <= MUX_s_1_2_2({exit_ACC1_for_lpi_2_dfm_1 , ((MUX_s_1_2_2({(~
            (ACC1_for_acc_itm[2])) , exit_ACC1_for_lpi_2_dfm_1}, or_dcpl_80 | (~
            FRAME_stage_0))) | (exit_SHIFT_lpi_2_dfm_2 & ACC1_for_nand_tmp & FRAME_stage_0))},
            fsm_output[1]);
        regs_operator_din_lpi_2 <= regs_operator_din_lpi_2_mx0;
        apply_lpi_2_dfm_2 <= apply_lpi_2_dfm_1;
        exit_SHIFT_lpi_2_dfm_1 <= exit_SHIFT_lpi_2_dfm_2;
        ACC1_for_j_1_lpi_2_dfm_4 <= ACC1_for_j_1_lpi_2_dfm_4_mx1w0;
        i_1_lpi_2_dfm_2 <= i_1_lpi_2_dfm_2_mx1w0;
        exit_ACC1_lpi_2_dfm_3 <= exit_ACC1_lpi_2_dfm_1_mx0;
        regs_regs_4_lpi_2_dfm_1 <= regs_regs_4_lpi_2;
        regs_regs_3_lpi_2_dfm_1 <= regs_regs_3_lpi_2;
        regs_regs_2_lpi_2_dfm_1 <= regs_regs_2_lpi_2;
        regs_regs_1_lpi_2_dfm_1 <= regs_regs_1_lpi_2;
        regs_regs_0_lpi_2_dfm_1 <= regs_regs_0_lpi_2;
      end
    end
  end

  function [2:0] MUX_v_3_2_2;
    input [5:0] inputs;
    input [0:0] sel;
    reg [2:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[5:3];
      end
      1'b1 : begin
        result = inputs[2:0];
      end
      default : begin
        result = inputs[5:3];
      end
    endcase
    MUX_v_3_2_2 = result;
  end
  endfunction


  function [2:0] signext_3_1;
    input [0:0] vector;
  begin
    signext_3_1= {{2{vector[0]}}, vector};
  end
  endfunction


  function [0:0] MUX_s_1_2_2;
    input [1:0] inputs;
    input [0:0] sel;
    reg [0:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[1:1];
      end
      1'b1 : begin
        result = inputs[0:0];
      end
      default : begin
        result = inputs[1:1];
      end
    endcase
    MUX_s_1_2_2 = result;
  end
  endfunction


  function [149:0] MUX_v_150_2_2;
    input [299:0] inputs;
    input [0:0] sel;
    reg [149:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[299:150];
      end
      1'b1 : begin
        result = inputs[149:0];
      end
      default : begin
        result = inputs[299:150];
      end
    endcase
    MUX_v_150_2_2 = result;
  end
  endfunction


  function [1:0] MUX_v_2_512_2;
    input [1023:0] inputs;
    input [8:0] sel;
    reg [1:0] result;
  begin
    case (sel)
      9'b000000000 : begin
        result = inputs[1023:1022];
      end
      9'b000000001 : begin
        result = inputs[1021:1020];
      end
      9'b000000010 : begin
        result = inputs[1019:1018];
      end
      9'b000000011 : begin
        result = inputs[1017:1016];
      end
      9'b000000100 : begin
        result = inputs[1015:1014];
      end
      9'b000000101 : begin
        result = inputs[1013:1012];
      end
      9'b000000110 : begin
        result = inputs[1011:1010];
      end
      9'b000000111 : begin
        result = inputs[1009:1008];
      end
      9'b000001000 : begin
        result = inputs[1007:1006];
      end
      9'b000001001 : begin
        result = inputs[1005:1004];
      end
      9'b000001010 : begin
        result = inputs[1003:1002];
      end
      9'b000001011 : begin
        result = inputs[1001:1000];
      end
      9'b000001100 : begin
        result = inputs[999:998];
      end
      9'b000001101 : begin
        result = inputs[997:996];
      end
      9'b000001110 : begin
        result = inputs[995:994];
      end
      9'b000001111 : begin
        result = inputs[993:992];
      end
      9'b000010000 : begin
        result = inputs[991:990];
      end
      9'b000010001 : begin
        result = inputs[989:988];
      end
      9'b000010010 : begin
        result = inputs[987:986];
      end
      9'b000010011 : begin
        result = inputs[985:984];
      end
      9'b000010100 : begin
        result = inputs[983:982];
      end
      9'b000010101 : begin
        result = inputs[981:980];
      end
      9'b000010110 : begin
        result = inputs[979:978];
      end
      9'b000010111 : begin
        result = inputs[977:976];
      end
      9'b000011000 : begin
        result = inputs[975:974];
      end
      9'b000011001 : begin
        result = inputs[973:972];
      end
      9'b000011010 : begin
        result = inputs[971:970];
      end
      9'b000011011 : begin
        result = inputs[969:968];
      end
      9'b000011100 : begin
        result = inputs[967:966];
      end
      9'b000011101 : begin
        result = inputs[965:964];
      end
      9'b000011110 : begin
        result = inputs[963:962];
      end
      9'b000011111 : begin
        result = inputs[961:960];
      end
      9'b000100000 : begin
        result = inputs[959:958];
      end
      9'b000100001 : begin
        result = inputs[957:956];
      end
      9'b000100010 : begin
        result = inputs[955:954];
      end
      9'b000100011 : begin
        result = inputs[953:952];
      end
      9'b000100100 : begin
        result = inputs[951:950];
      end
      9'b000100101 : begin
        result = inputs[949:948];
      end
      9'b000100110 : begin
        result = inputs[947:946];
      end
      9'b000100111 : begin
        result = inputs[945:944];
      end
      9'b000101000 : begin
        result = inputs[943:942];
      end
      9'b000101001 : begin
        result = inputs[941:940];
      end
      9'b000101010 : begin
        result = inputs[939:938];
      end
      9'b000101011 : begin
        result = inputs[937:936];
      end
      9'b000101100 : begin
        result = inputs[935:934];
      end
      9'b000101101 : begin
        result = inputs[933:932];
      end
      9'b000101110 : begin
        result = inputs[931:930];
      end
      9'b000101111 : begin
        result = inputs[929:928];
      end
      9'b000110000 : begin
        result = inputs[927:926];
      end
      9'b000110001 : begin
        result = inputs[925:924];
      end
      9'b000110010 : begin
        result = inputs[923:922];
      end
      9'b000110011 : begin
        result = inputs[921:920];
      end
      9'b000110100 : begin
        result = inputs[919:918];
      end
      9'b000110101 : begin
        result = inputs[917:916];
      end
      9'b000110110 : begin
        result = inputs[915:914];
      end
      9'b000110111 : begin
        result = inputs[913:912];
      end
      9'b000111000 : begin
        result = inputs[911:910];
      end
      9'b000111001 : begin
        result = inputs[909:908];
      end
      9'b000111010 : begin
        result = inputs[907:906];
      end
      9'b000111011 : begin
        result = inputs[905:904];
      end
      9'b000111100 : begin
        result = inputs[903:902];
      end
      9'b000111101 : begin
        result = inputs[901:900];
      end
      9'b000111110 : begin
        result = inputs[899:898];
      end
      9'b000111111 : begin
        result = inputs[897:896];
      end
      9'b001000000 : begin
        result = inputs[895:894];
      end
      9'b001000001 : begin
        result = inputs[893:892];
      end
      9'b001000010 : begin
        result = inputs[891:890];
      end
      9'b001000011 : begin
        result = inputs[889:888];
      end
      9'b001000100 : begin
        result = inputs[887:886];
      end
      9'b001000101 : begin
        result = inputs[885:884];
      end
      9'b001000110 : begin
        result = inputs[883:882];
      end
      9'b001000111 : begin
        result = inputs[881:880];
      end
      9'b001001000 : begin
        result = inputs[879:878];
      end
      9'b001001001 : begin
        result = inputs[877:876];
      end
      9'b001001010 : begin
        result = inputs[875:874];
      end
      9'b001001011 : begin
        result = inputs[873:872];
      end
      9'b001001100 : begin
        result = inputs[871:870];
      end
      9'b001001101 : begin
        result = inputs[869:868];
      end
      9'b001001110 : begin
        result = inputs[867:866];
      end
      9'b001001111 : begin
        result = inputs[865:864];
      end
      9'b001010000 : begin
        result = inputs[863:862];
      end
      9'b001010001 : begin
        result = inputs[861:860];
      end
      9'b001010010 : begin
        result = inputs[859:858];
      end
      9'b001010011 : begin
        result = inputs[857:856];
      end
      9'b001010100 : begin
        result = inputs[855:854];
      end
      9'b001010101 : begin
        result = inputs[853:852];
      end
      9'b001010110 : begin
        result = inputs[851:850];
      end
      9'b001010111 : begin
        result = inputs[849:848];
      end
      9'b001011000 : begin
        result = inputs[847:846];
      end
      9'b001011001 : begin
        result = inputs[845:844];
      end
      9'b001011010 : begin
        result = inputs[843:842];
      end
      9'b001011011 : begin
        result = inputs[841:840];
      end
      9'b001011100 : begin
        result = inputs[839:838];
      end
      9'b001011101 : begin
        result = inputs[837:836];
      end
      9'b001011110 : begin
        result = inputs[835:834];
      end
      9'b001011111 : begin
        result = inputs[833:832];
      end
      9'b001100000 : begin
        result = inputs[831:830];
      end
      9'b001100001 : begin
        result = inputs[829:828];
      end
      9'b001100010 : begin
        result = inputs[827:826];
      end
      9'b001100011 : begin
        result = inputs[825:824];
      end
      9'b001100100 : begin
        result = inputs[823:822];
      end
      9'b001100101 : begin
        result = inputs[821:820];
      end
      9'b001100110 : begin
        result = inputs[819:818];
      end
      9'b001100111 : begin
        result = inputs[817:816];
      end
      9'b001101000 : begin
        result = inputs[815:814];
      end
      9'b001101001 : begin
        result = inputs[813:812];
      end
      9'b001101010 : begin
        result = inputs[811:810];
      end
      9'b001101011 : begin
        result = inputs[809:808];
      end
      9'b001101100 : begin
        result = inputs[807:806];
      end
      9'b001101101 : begin
        result = inputs[805:804];
      end
      9'b001101110 : begin
        result = inputs[803:802];
      end
      9'b001101111 : begin
        result = inputs[801:800];
      end
      9'b001110000 : begin
        result = inputs[799:798];
      end
      9'b001110001 : begin
        result = inputs[797:796];
      end
      9'b001110010 : begin
        result = inputs[795:794];
      end
      9'b001110011 : begin
        result = inputs[793:792];
      end
      9'b001110100 : begin
        result = inputs[791:790];
      end
      9'b001110101 : begin
        result = inputs[789:788];
      end
      9'b001110110 : begin
        result = inputs[787:786];
      end
      9'b001110111 : begin
        result = inputs[785:784];
      end
      9'b001111000 : begin
        result = inputs[783:782];
      end
      9'b001111001 : begin
        result = inputs[781:780];
      end
      9'b001111010 : begin
        result = inputs[779:778];
      end
      9'b001111011 : begin
        result = inputs[777:776];
      end
      9'b001111100 : begin
        result = inputs[775:774];
      end
      9'b001111101 : begin
        result = inputs[773:772];
      end
      9'b001111110 : begin
        result = inputs[771:770];
      end
      9'b001111111 : begin
        result = inputs[769:768];
      end
      9'b010000000 : begin
        result = inputs[767:766];
      end
      9'b010000001 : begin
        result = inputs[765:764];
      end
      9'b010000010 : begin
        result = inputs[763:762];
      end
      9'b010000011 : begin
        result = inputs[761:760];
      end
      9'b010000100 : begin
        result = inputs[759:758];
      end
      9'b010000101 : begin
        result = inputs[757:756];
      end
      9'b010000110 : begin
        result = inputs[755:754];
      end
      9'b010000111 : begin
        result = inputs[753:752];
      end
      9'b010001000 : begin
        result = inputs[751:750];
      end
      9'b010001001 : begin
        result = inputs[749:748];
      end
      9'b010001010 : begin
        result = inputs[747:746];
      end
      9'b010001011 : begin
        result = inputs[745:744];
      end
      9'b010001100 : begin
        result = inputs[743:742];
      end
      9'b010001101 : begin
        result = inputs[741:740];
      end
      9'b010001110 : begin
        result = inputs[739:738];
      end
      9'b010001111 : begin
        result = inputs[737:736];
      end
      9'b010010000 : begin
        result = inputs[735:734];
      end
      9'b010010001 : begin
        result = inputs[733:732];
      end
      9'b010010010 : begin
        result = inputs[731:730];
      end
      9'b010010011 : begin
        result = inputs[729:728];
      end
      9'b010010100 : begin
        result = inputs[727:726];
      end
      9'b010010101 : begin
        result = inputs[725:724];
      end
      9'b010010110 : begin
        result = inputs[723:722];
      end
      9'b010010111 : begin
        result = inputs[721:720];
      end
      9'b010011000 : begin
        result = inputs[719:718];
      end
      9'b010011001 : begin
        result = inputs[717:716];
      end
      9'b010011010 : begin
        result = inputs[715:714];
      end
      9'b010011011 : begin
        result = inputs[713:712];
      end
      9'b010011100 : begin
        result = inputs[711:710];
      end
      9'b010011101 : begin
        result = inputs[709:708];
      end
      9'b010011110 : begin
        result = inputs[707:706];
      end
      9'b010011111 : begin
        result = inputs[705:704];
      end
      9'b010100000 : begin
        result = inputs[703:702];
      end
      9'b010100001 : begin
        result = inputs[701:700];
      end
      9'b010100010 : begin
        result = inputs[699:698];
      end
      9'b010100011 : begin
        result = inputs[697:696];
      end
      9'b010100100 : begin
        result = inputs[695:694];
      end
      9'b010100101 : begin
        result = inputs[693:692];
      end
      9'b010100110 : begin
        result = inputs[691:690];
      end
      9'b010100111 : begin
        result = inputs[689:688];
      end
      9'b010101000 : begin
        result = inputs[687:686];
      end
      9'b010101001 : begin
        result = inputs[685:684];
      end
      9'b010101010 : begin
        result = inputs[683:682];
      end
      9'b010101011 : begin
        result = inputs[681:680];
      end
      9'b010101100 : begin
        result = inputs[679:678];
      end
      9'b010101101 : begin
        result = inputs[677:676];
      end
      9'b010101110 : begin
        result = inputs[675:674];
      end
      9'b010101111 : begin
        result = inputs[673:672];
      end
      9'b010110000 : begin
        result = inputs[671:670];
      end
      9'b010110001 : begin
        result = inputs[669:668];
      end
      9'b010110010 : begin
        result = inputs[667:666];
      end
      9'b010110011 : begin
        result = inputs[665:664];
      end
      9'b010110100 : begin
        result = inputs[663:662];
      end
      9'b010110101 : begin
        result = inputs[661:660];
      end
      9'b010110110 : begin
        result = inputs[659:658];
      end
      9'b010110111 : begin
        result = inputs[657:656];
      end
      9'b010111000 : begin
        result = inputs[655:654];
      end
      9'b010111001 : begin
        result = inputs[653:652];
      end
      9'b010111010 : begin
        result = inputs[651:650];
      end
      9'b010111011 : begin
        result = inputs[649:648];
      end
      9'b010111100 : begin
        result = inputs[647:646];
      end
      9'b010111101 : begin
        result = inputs[645:644];
      end
      9'b010111110 : begin
        result = inputs[643:642];
      end
      9'b010111111 : begin
        result = inputs[641:640];
      end
      9'b011000000 : begin
        result = inputs[639:638];
      end
      9'b011000001 : begin
        result = inputs[637:636];
      end
      9'b011000010 : begin
        result = inputs[635:634];
      end
      9'b011000011 : begin
        result = inputs[633:632];
      end
      9'b011000100 : begin
        result = inputs[631:630];
      end
      9'b011000101 : begin
        result = inputs[629:628];
      end
      9'b011000110 : begin
        result = inputs[627:626];
      end
      9'b011000111 : begin
        result = inputs[625:624];
      end
      9'b011001000 : begin
        result = inputs[623:622];
      end
      9'b011001001 : begin
        result = inputs[621:620];
      end
      9'b011001010 : begin
        result = inputs[619:618];
      end
      9'b011001011 : begin
        result = inputs[617:616];
      end
      9'b011001100 : begin
        result = inputs[615:614];
      end
      9'b011001101 : begin
        result = inputs[613:612];
      end
      9'b011001110 : begin
        result = inputs[611:610];
      end
      9'b011001111 : begin
        result = inputs[609:608];
      end
      9'b011010000 : begin
        result = inputs[607:606];
      end
      9'b011010001 : begin
        result = inputs[605:604];
      end
      9'b011010010 : begin
        result = inputs[603:602];
      end
      9'b011010011 : begin
        result = inputs[601:600];
      end
      9'b011010100 : begin
        result = inputs[599:598];
      end
      9'b011010101 : begin
        result = inputs[597:596];
      end
      9'b011010110 : begin
        result = inputs[595:594];
      end
      9'b011010111 : begin
        result = inputs[593:592];
      end
      9'b011011000 : begin
        result = inputs[591:590];
      end
      9'b011011001 : begin
        result = inputs[589:588];
      end
      9'b011011010 : begin
        result = inputs[587:586];
      end
      9'b011011011 : begin
        result = inputs[585:584];
      end
      9'b011011100 : begin
        result = inputs[583:582];
      end
      9'b011011101 : begin
        result = inputs[581:580];
      end
      9'b011011110 : begin
        result = inputs[579:578];
      end
      9'b011011111 : begin
        result = inputs[577:576];
      end
      9'b011100000 : begin
        result = inputs[575:574];
      end
      9'b011100001 : begin
        result = inputs[573:572];
      end
      9'b011100010 : begin
        result = inputs[571:570];
      end
      9'b011100011 : begin
        result = inputs[569:568];
      end
      9'b011100100 : begin
        result = inputs[567:566];
      end
      9'b011100101 : begin
        result = inputs[565:564];
      end
      9'b011100110 : begin
        result = inputs[563:562];
      end
      9'b011100111 : begin
        result = inputs[561:560];
      end
      9'b011101000 : begin
        result = inputs[559:558];
      end
      9'b011101001 : begin
        result = inputs[557:556];
      end
      9'b011101010 : begin
        result = inputs[555:554];
      end
      9'b011101011 : begin
        result = inputs[553:552];
      end
      9'b011101100 : begin
        result = inputs[551:550];
      end
      9'b011101101 : begin
        result = inputs[549:548];
      end
      9'b011101110 : begin
        result = inputs[547:546];
      end
      9'b011101111 : begin
        result = inputs[545:544];
      end
      9'b011110000 : begin
        result = inputs[543:542];
      end
      9'b011110001 : begin
        result = inputs[541:540];
      end
      9'b011110010 : begin
        result = inputs[539:538];
      end
      9'b011110011 : begin
        result = inputs[537:536];
      end
      9'b011110100 : begin
        result = inputs[535:534];
      end
      9'b011110101 : begin
        result = inputs[533:532];
      end
      9'b011110110 : begin
        result = inputs[531:530];
      end
      9'b011110111 : begin
        result = inputs[529:528];
      end
      9'b011111000 : begin
        result = inputs[527:526];
      end
      9'b011111001 : begin
        result = inputs[525:524];
      end
      9'b011111010 : begin
        result = inputs[523:522];
      end
      9'b011111011 : begin
        result = inputs[521:520];
      end
      9'b011111100 : begin
        result = inputs[519:518];
      end
      9'b011111101 : begin
        result = inputs[517:516];
      end
      9'b011111110 : begin
        result = inputs[515:514];
      end
      9'b011111111 : begin
        result = inputs[513:512];
      end
      9'b100000000 : begin
        result = inputs[511:510];
      end
      9'b100000001 : begin
        result = inputs[509:508];
      end
      9'b100000010 : begin
        result = inputs[507:506];
      end
      9'b100000011 : begin
        result = inputs[505:504];
      end
      9'b100000100 : begin
        result = inputs[503:502];
      end
      9'b100000101 : begin
        result = inputs[501:500];
      end
      9'b100000110 : begin
        result = inputs[499:498];
      end
      9'b100000111 : begin
        result = inputs[497:496];
      end
      9'b100001000 : begin
        result = inputs[495:494];
      end
      9'b100001001 : begin
        result = inputs[493:492];
      end
      9'b100001010 : begin
        result = inputs[491:490];
      end
      9'b100001011 : begin
        result = inputs[489:488];
      end
      9'b100001100 : begin
        result = inputs[487:486];
      end
      9'b100001101 : begin
        result = inputs[485:484];
      end
      9'b100001110 : begin
        result = inputs[483:482];
      end
      9'b100001111 : begin
        result = inputs[481:480];
      end
      9'b100010000 : begin
        result = inputs[479:478];
      end
      9'b100010001 : begin
        result = inputs[477:476];
      end
      9'b100010010 : begin
        result = inputs[475:474];
      end
      9'b100010011 : begin
        result = inputs[473:472];
      end
      9'b100010100 : begin
        result = inputs[471:470];
      end
      9'b100010101 : begin
        result = inputs[469:468];
      end
      9'b100010110 : begin
        result = inputs[467:466];
      end
      9'b100010111 : begin
        result = inputs[465:464];
      end
      9'b100011000 : begin
        result = inputs[463:462];
      end
      9'b100011001 : begin
        result = inputs[461:460];
      end
      9'b100011010 : begin
        result = inputs[459:458];
      end
      9'b100011011 : begin
        result = inputs[457:456];
      end
      9'b100011100 : begin
        result = inputs[455:454];
      end
      9'b100011101 : begin
        result = inputs[453:452];
      end
      9'b100011110 : begin
        result = inputs[451:450];
      end
      9'b100011111 : begin
        result = inputs[449:448];
      end
      9'b100100000 : begin
        result = inputs[447:446];
      end
      9'b100100001 : begin
        result = inputs[445:444];
      end
      9'b100100010 : begin
        result = inputs[443:442];
      end
      9'b100100011 : begin
        result = inputs[441:440];
      end
      9'b100100100 : begin
        result = inputs[439:438];
      end
      9'b100100101 : begin
        result = inputs[437:436];
      end
      9'b100100110 : begin
        result = inputs[435:434];
      end
      9'b100100111 : begin
        result = inputs[433:432];
      end
      9'b100101000 : begin
        result = inputs[431:430];
      end
      9'b100101001 : begin
        result = inputs[429:428];
      end
      9'b100101010 : begin
        result = inputs[427:426];
      end
      9'b100101011 : begin
        result = inputs[425:424];
      end
      9'b100101100 : begin
        result = inputs[423:422];
      end
      9'b100101101 : begin
        result = inputs[421:420];
      end
      9'b100101110 : begin
        result = inputs[419:418];
      end
      9'b100101111 : begin
        result = inputs[417:416];
      end
      9'b100110000 : begin
        result = inputs[415:414];
      end
      9'b100110001 : begin
        result = inputs[413:412];
      end
      9'b100110010 : begin
        result = inputs[411:410];
      end
      9'b100110011 : begin
        result = inputs[409:408];
      end
      9'b100110100 : begin
        result = inputs[407:406];
      end
      9'b100110101 : begin
        result = inputs[405:404];
      end
      9'b100110110 : begin
        result = inputs[403:402];
      end
      9'b100110111 : begin
        result = inputs[401:400];
      end
      9'b100111000 : begin
        result = inputs[399:398];
      end
      9'b100111001 : begin
        result = inputs[397:396];
      end
      9'b100111010 : begin
        result = inputs[395:394];
      end
      9'b100111011 : begin
        result = inputs[393:392];
      end
      9'b100111100 : begin
        result = inputs[391:390];
      end
      9'b100111101 : begin
        result = inputs[389:388];
      end
      9'b100111110 : begin
        result = inputs[387:386];
      end
      9'b100111111 : begin
        result = inputs[385:384];
      end
      9'b101000000 : begin
        result = inputs[383:382];
      end
      9'b101000001 : begin
        result = inputs[381:380];
      end
      9'b101000010 : begin
        result = inputs[379:378];
      end
      9'b101000011 : begin
        result = inputs[377:376];
      end
      9'b101000100 : begin
        result = inputs[375:374];
      end
      9'b101000101 : begin
        result = inputs[373:372];
      end
      9'b101000110 : begin
        result = inputs[371:370];
      end
      9'b101000111 : begin
        result = inputs[369:368];
      end
      9'b101001000 : begin
        result = inputs[367:366];
      end
      9'b101001001 : begin
        result = inputs[365:364];
      end
      9'b101001010 : begin
        result = inputs[363:362];
      end
      9'b101001011 : begin
        result = inputs[361:360];
      end
      9'b101001100 : begin
        result = inputs[359:358];
      end
      9'b101001101 : begin
        result = inputs[357:356];
      end
      9'b101001110 : begin
        result = inputs[355:354];
      end
      9'b101001111 : begin
        result = inputs[353:352];
      end
      9'b101010000 : begin
        result = inputs[351:350];
      end
      9'b101010001 : begin
        result = inputs[349:348];
      end
      9'b101010010 : begin
        result = inputs[347:346];
      end
      9'b101010011 : begin
        result = inputs[345:344];
      end
      9'b101010100 : begin
        result = inputs[343:342];
      end
      9'b101010101 : begin
        result = inputs[341:340];
      end
      9'b101010110 : begin
        result = inputs[339:338];
      end
      9'b101010111 : begin
        result = inputs[337:336];
      end
      9'b101011000 : begin
        result = inputs[335:334];
      end
      9'b101011001 : begin
        result = inputs[333:332];
      end
      9'b101011010 : begin
        result = inputs[331:330];
      end
      9'b101011011 : begin
        result = inputs[329:328];
      end
      9'b101011100 : begin
        result = inputs[327:326];
      end
      9'b101011101 : begin
        result = inputs[325:324];
      end
      9'b101011110 : begin
        result = inputs[323:322];
      end
      9'b101011111 : begin
        result = inputs[321:320];
      end
      9'b101100000 : begin
        result = inputs[319:318];
      end
      9'b101100001 : begin
        result = inputs[317:316];
      end
      9'b101100010 : begin
        result = inputs[315:314];
      end
      9'b101100011 : begin
        result = inputs[313:312];
      end
      9'b101100100 : begin
        result = inputs[311:310];
      end
      9'b101100101 : begin
        result = inputs[309:308];
      end
      9'b101100110 : begin
        result = inputs[307:306];
      end
      9'b101100111 : begin
        result = inputs[305:304];
      end
      9'b101101000 : begin
        result = inputs[303:302];
      end
      9'b101101001 : begin
        result = inputs[301:300];
      end
      9'b101101010 : begin
        result = inputs[299:298];
      end
      9'b101101011 : begin
        result = inputs[297:296];
      end
      9'b101101100 : begin
        result = inputs[295:294];
      end
      9'b101101101 : begin
        result = inputs[293:292];
      end
      9'b101101110 : begin
        result = inputs[291:290];
      end
      9'b101101111 : begin
        result = inputs[289:288];
      end
      9'b101110000 : begin
        result = inputs[287:286];
      end
      9'b101110001 : begin
        result = inputs[285:284];
      end
      9'b101110010 : begin
        result = inputs[283:282];
      end
      9'b101110011 : begin
        result = inputs[281:280];
      end
      9'b101110100 : begin
        result = inputs[279:278];
      end
      9'b101110101 : begin
        result = inputs[277:276];
      end
      9'b101110110 : begin
        result = inputs[275:274];
      end
      9'b101110111 : begin
        result = inputs[273:272];
      end
      9'b101111000 : begin
        result = inputs[271:270];
      end
      9'b101111001 : begin
        result = inputs[269:268];
      end
      9'b101111010 : begin
        result = inputs[267:266];
      end
      9'b101111011 : begin
        result = inputs[265:264];
      end
      9'b101111100 : begin
        result = inputs[263:262];
      end
      9'b101111101 : begin
        result = inputs[261:260];
      end
      9'b101111110 : begin
        result = inputs[259:258];
      end
      9'b101111111 : begin
        result = inputs[257:256];
      end
      9'b110000000 : begin
        result = inputs[255:254];
      end
      9'b110000001 : begin
        result = inputs[253:252];
      end
      9'b110000010 : begin
        result = inputs[251:250];
      end
      9'b110000011 : begin
        result = inputs[249:248];
      end
      9'b110000100 : begin
        result = inputs[247:246];
      end
      9'b110000101 : begin
        result = inputs[245:244];
      end
      9'b110000110 : begin
        result = inputs[243:242];
      end
      9'b110000111 : begin
        result = inputs[241:240];
      end
      9'b110001000 : begin
        result = inputs[239:238];
      end
      9'b110001001 : begin
        result = inputs[237:236];
      end
      9'b110001010 : begin
        result = inputs[235:234];
      end
      9'b110001011 : begin
        result = inputs[233:232];
      end
      9'b110001100 : begin
        result = inputs[231:230];
      end
      9'b110001101 : begin
        result = inputs[229:228];
      end
      9'b110001110 : begin
        result = inputs[227:226];
      end
      9'b110001111 : begin
        result = inputs[225:224];
      end
      9'b110010000 : begin
        result = inputs[223:222];
      end
      9'b110010001 : begin
        result = inputs[221:220];
      end
      9'b110010010 : begin
        result = inputs[219:218];
      end
      9'b110010011 : begin
        result = inputs[217:216];
      end
      9'b110010100 : begin
        result = inputs[215:214];
      end
      9'b110010101 : begin
        result = inputs[213:212];
      end
      9'b110010110 : begin
        result = inputs[211:210];
      end
      9'b110010111 : begin
        result = inputs[209:208];
      end
      9'b110011000 : begin
        result = inputs[207:206];
      end
      9'b110011001 : begin
        result = inputs[205:204];
      end
      9'b110011010 : begin
        result = inputs[203:202];
      end
      9'b110011011 : begin
        result = inputs[201:200];
      end
      9'b110011100 : begin
        result = inputs[199:198];
      end
      9'b110011101 : begin
        result = inputs[197:196];
      end
      9'b110011110 : begin
        result = inputs[195:194];
      end
      9'b110011111 : begin
        result = inputs[193:192];
      end
      9'b110100000 : begin
        result = inputs[191:190];
      end
      9'b110100001 : begin
        result = inputs[189:188];
      end
      9'b110100010 : begin
        result = inputs[187:186];
      end
      9'b110100011 : begin
        result = inputs[185:184];
      end
      9'b110100100 : begin
        result = inputs[183:182];
      end
      9'b110100101 : begin
        result = inputs[181:180];
      end
      9'b110100110 : begin
        result = inputs[179:178];
      end
      9'b110100111 : begin
        result = inputs[177:176];
      end
      9'b110101000 : begin
        result = inputs[175:174];
      end
      9'b110101001 : begin
        result = inputs[173:172];
      end
      9'b110101010 : begin
        result = inputs[171:170];
      end
      9'b110101011 : begin
        result = inputs[169:168];
      end
      9'b110101100 : begin
        result = inputs[167:166];
      end
      9'b110101101 : begin
        result = inputs[165:164];
      end
      9'b110101110 : begin
        result = inputs[163:162];
      end
      9'b110101111 : begin
        result = inputs[161:160];
      end
      9'b110110000 : begin
        result = inputs[159:158];
      end
      9'b110110001 : begin
        result = inputs[157:156];
      end
      9'b110110010 : begin
        result = inputs[155:154];
      end
      9'b110110011 : begin
        result = inputs[153:152];
      end
      9'b110110100 : begin
        result = inputs[151:150];
      end
      9'b110110101 : begin
        result = inputs[149:148];
      end
      9'b110110110 : begin
        result = inputs[147:146];
      end
      9'b110110111 : begin
        result = inputs[145:144];
      end
      9'b110111000 : begin
        result = inputs[143:142];
      end
      9'b110111001 : begin
        result = inputs[141:140];
      end
      9'b110111010 : begin
        result = inputs[139:138];
      end
      9'b110111011 : begin
        result = inputs[137:136];
      end
      9'b110111100 : begin
        result = inputs[135:134];
      end
      9'b110111101 : begin
        result = inputs[133:132];
      end
      9'b110111110 : begin
        result = inputs[131:130];
      end
      9'b110111111 : begin
        result = inputs[129:128];
      end
      9'b111000000 : begin
        result = inputs[127:126];
      end
      9'b111000001 : begin
        result = inputs[125:124];
      end
      9'b111000010 : begin
        result = inputs[123:122];
      end
      9'b111000011 : begin
        result = inputs[121:120];
      end
      9'b111000100 : begin
        result = inputs[119:118];
      end
      9'b111000101 : begin
        result = inputs[117:116];
      end
      9'b111000110 : begin
        result = inputs[115:114];
      end
      9'b111000111 : begin
        result = inputs[113:112];
      end
      9'b111001000 : begin
        result = inputs[111:110];
      end
      9'b111001001 : begin
        result = inputs[109:108];
      end
      9'b111001010 : begin
        result = inputs[107:106];
      end
      9'b111001011 : begin
        result = inputs[105:104];
      end
      9'b111001100 : begin
        result = inputs[103:102];
      end
      9'b111001101 : begin
        result = inputs[101:100];
      end
      9'b111001110 : begin
        result = inputs[99:98];
      end
      9'b111001111 : begin
        result = inputs[97:96];
      end
      9'b111010000 : begin
        result = inputs[95:94];
      end
      9'b111010001 : begin
        result = inputs[93:92];
      end
      9'b111010010 : begin
        result = inputs[91:90];
      end
      9'b111010011 : begin
        result = inputs[89:88];
      end
      9'b111010100 : begin
        result = inputs[87:86];
      end
      9'b111010101 : begin
        result = inputs[85:84];
      end
      9'b111010110 : begin
        result = inputs[83:82];
      end
      9'b111010111 : begin
        result = inputs[81:80];
      end
      9'b111011000 : begin
        result = inputs[79:78];
      end
      9'b111011001 : begin
        result = inputs[77:76];
      end
      9'b111011010 : begin
        result = inputs[75:74];
      end
      9'b111011011 : begin
        result = inputs[73:72];
      end
      9'b111011100 : begin
        result = inputs[71:70];
      end
      9'b111011101 : begin
        result = inputs[69:68];
      end
      9'b111011110 : begin
        result = inputs[67:66];
      end
      9'b111011111 : begin
        result = inputs[65:64];
      end
      9'b111100000 : begin
        result = inputs[63:62];
      end
      9'b111100001 : begin
        result = inputs[61:60];
      end
      9'b111100010 : begin
        result = inputs[59:58];
      end
      9'b111100011 : begin
        result = inputs[57:56];
      end
      9'b111100100 : begin
        result = inputs[55:54];
      end
      9'b111100101 : begin
        result = inputs[53:52];
      end
      9'b111100110 : begin
        result = inputs[51:50];
      end
      9'b111100111 : begin
        result = inputs[49:48];
      end
      9'b111101000 : begin
        result = inputs[47:46];
      end
      9'b111101001 : begin
        result = inputs[45:44];
      end
      9'b111101010 : begin
        result = inputs[43:42];
      end
      9'b111101011 : begin
        result = inputs[41:40];
      end
      9'b111101100 : begin
        result = inputs[39:38];
      end
      9'b111101101 : begin
        result = inputs[37:36];
      end
      9'b111101110 : begin
        result = inputs[35:34];
      end
      9'b111101111 : begin
        result = inputs[33:32];
      end
      9'b111110000 : begin
        result = inputs[31:30];
      end
      9'b111110001 : begin
        result = inputs[29:28];
      end
      9'b111110010 : begin
        result = inputs[27:26];
      end
      9'b111110011 : begin
        result = inputs[25:24];
      end
      9'b111110100 : begin
        result = inputs[23:22];
      end
      9'b111110101 : begin
        result = inputs[21:20];
      end
      9'b111110110 : begin
        result = inputs[19:18];
      end
      9'b111110111 : begin
        result = inputs[17:16];
      end
      9'b111111000 : begin
        result = inputs[15:14];
      end
      9'b111111001 : begin
        result = inputs[13:12];
      end
      9'b111111010 : begin
        result = inputs[11:10];
      end
      9'b111111011 : begin
        result = inputs[9:8];
      end
      9'b111111100 : begin
        result = inputs[7:6];
      end
      9'b111111101 : begin
        result = inputs[5:4];
      end
      9'b111111110 : begin
        result = inputs[3:2];
      end
      9'b111111111 : begin
        result = inputs[1:0];
      end
      default : begin
        result = inputs[1023:1022];
      end
    endcase
    MUX_v_2_512_2 = result;
  end
  endfunction


  function [149:0] MUX_v_150_4_2;
    input [599:0] inputs;
    input [1:0] sel;
    reg [149:0] result;
  begin
    case (sel)
      2'b00 : begin
        result = inputs[599:450];
      end
      2'b01 : begin
        result = inputs[449:300];
      end
      2'b10 : begin
        result = inputs[299:150];
      end
      2'b11 : begin
        result = inputs[149:0];
      end
      default : begin
        result = inputs[599:450];
      end
    endcase
    MUX_v_150_4_2 = result;
  end
  endfunction


  function [29:0] signext_30_1;
    input [0:0] vector;
  begin
    signext_30_1= {{29{vector[0]}}, vector};
  end
  endfunction


  function [0:0] readslicef_8_1_7;
    input [7:0] vector;
    reg [7:0] tmp;
  begin
    tmp = vector >> 7;
    readslicef_8_1_7 = tmp[0:0];
  end
  endfunction


  function [18:0] MUX_v_19_2_2;
    input [37:0] inputs;
    input [0:0] sel;
    reg [18:0] result;
  begin
    case (sel)
      1'b0 : begin
        result = inputs[37:19];
      end
      1'b1 : begin
        result = inputs[18:0];
      end
      default : begin
        result = inputs[37:19];
      end
    endcase
    MUX_v_19_2_2 = result;
  end
  endfunction


  function [18:0] signext_19_1;
    input [0:0] vector;
  begin
    signext_19_1= {{18{vector[0]}}, vector};
  end
  endfunction


  function [2:0] MUX1HOT_v_3_3_2;
    input [8:0] inputs;
    input [2:0] sel;
    reg [2:0] result;
    integer i;
  begin
    result = inputs[0+:3] & {3{sel[0]}};
    for( i = 1; i < 3; i = i + 1 )
      result = result | (inputs[i*3+:3] & {3{sel[i]}});
    MUX1HOT_v_3_3_2 = result;
  end
  endfunction


  function [0:0] MUX1HOT_s_1_3_2;
    input [2:0] inputs;
    input [2:0] sel;
    reg [0:0] result;
    integer i;
  begin
    result = inputs[0+:1] & {1{sel[0]}};
    for( i = 1; i < 3; i = i + 1 )
      result = result | (inputs[i*1+:1] & {1{sel[i]}});
    MUX1HOT_s_1_3_2 = result;
  end
  endfunction


  function [149:0] MUX1HOT_v_150_3_2;
    input [449:0] inputs;
    input [2:0] sel;
    reg [149:0] result;
    integer i;
  begin
    result = inputs[0+:150] & {150{sel[0]}};
    for( i = 1; i < 3; i = i + 1 )
      result = result | (inputs[i*150+:150] & {150{sel[i]}});
    MUX1HOT_v_150_3_2 = result;
  end
  endfunction


  function  [8:0] conv_u2u_6_9 ;
    input [5:0]  vector ;
  begin
    conv_u2u_6_9 = {{3{1'b0}}, vector};
  end
  endfunction


  function  [5:0] conv_s2u_4_6 ;
    input signed [3:0]  vector ;
  begin
    conv_s2u_4_6 = {{2{vector[3]}}, vector};
  end
  endfunction


  function  [8:0] conv_u2u_18_9 ;
    input [17:0]  vector ;
  begin
    conv_u2u_18_9 = vector[8:0];
  end
  endfunction


  function  [8:0] conv_u2u_3_9 ;
    input [2:0]  vector ;
  begin
    conv_u2u_3_9 = {{6{1'b0}}, vector};
  end
  endfunction


  function signed [7:0] conv_u2s_7_8 ;
    input [6:0]  vector ;
  begin
    conv_u2s_7_8 = {1'b0, vector};
  end
  endfunction

endmodule

// ------------------------------------------------------------------
//  Design Unit:    erosion
//  Generated from file(s):
//    3) $PROJECT_HOME/erosion.c
// ------------------------------------------------------------------


module erosion (
  vin_rsc_z, vout_rsc_z, clk, en, arst_n
);
  input [149:0] vin_rsc_z;
  output [29:0] vout_rsc_z;
  input clk;
  input en;
  input arst_n;


  // Interconnect Declarations
  wire [149:0] vin_rsc_mgc_in_wire_d;
  wire [29:0] vout_rsc_mgc_out_stdreg_d;


  // Interconnect Declarations for Component Instantiations 
  mgc_in_wire #(.rscid(1),
  .width(150)) vin_rsc_mgc_in_wire (
      .d(vin_rsc_mgc_in_wire_d),
      .z(vin_rsc_z)
    );
  mgc_out_stdreg #(.rscid(2),
  .width(30)) vout_rsc_mgc_out_stdreg (
      .d(vout_rsc_mgc_out_stdreg_d),
      .z(vout_rsc_z)
    );
  erosion_core erosion_core_inst (
      .clk(clk),
      .en(en),
      .arst_n(arst_n),
      .vin_rsc_mgc_in_wire_d(vin_rsc_mgc_in_wire_d),
      .vout_rsc_mgc_out_stdreg_d(vout_rsc_mgc_out_stdreg_d)
    );
endmodule



